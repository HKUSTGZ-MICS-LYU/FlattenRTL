module top
    (
        input clk,
        input rst,
        input [127:0] state,
        input [127:0] key,
        output [127:0] out,
        output [63:0] Capacitance
    );
    wire \AES.clk ;
    wire [127:0] \AES.state ;
    wire [127:0] \AES.key ;
    wire [127:0] \AES.out ;
    reg [127:0] \AES.s0 ;
    reg [127:0] \AES.k0 ;
    wire [127:0] \AES.s1 ;
    wire [127:0] \AES.s2 ;
    wire [127:0] \AES.s3 ;
    wire [127:0] \AES.s4 ;
    wire [127:0] \AES.s5 ;
    wire [127:0] \AES.s6 ;
    wire [127:0] \AES.s7 ;
    wire [127:0] \AES.s8 ;
    wire [127:0] \AES.s9 ;
    wire [127:0] \AES.k1 ;
    wire [127:0] \AES.k2 ;
    wire [127:0] \AES.k3 ;
    wire [127:0] \AES.k4 ;
    wire [127:0] \AES.k5 ;
    wire [127:0] \AES.k6 ;
    wire [127:0] \AES.k7 ;
    wire [127:0] \AES.k8 ;
    wire [127:0] \AES.k9 ;
    wire [127:0] \AES.k10 ;
    wire [127:0] \AES.k0b ;
    wire [127:0] \AES.k1b ;
    wire [127:0] \AES.k2b ;
    wire [127:0] \AES.k3b ;
    wire [127:0] \AES.k4b ;
    wire [127:0] \AES.k5b ;
    wire [127:0] \AES.k6b ;
    wire [127:0] \AES.k7b ;
    wire [127:0] \AES.k8b ;
    wire [127:0] \AES.k9b ;
    wire [7:0] \AES.a1_rcon  = 8'h1;
    wire [7:0] \AES.a2_rcon  = 8'h2;
    wire [7:0] \AES.a3_rcon  = 8'h4;
    wire [7:0] \AES.a4_rcon  = 8'h8;
    wire [7:0] \AES.a5_rcon  = 8'h10;
    wire [7:0] \AES.a6_rcon  = 8'h20;
    wire [7:0] \AES.a7_rcon  = 8'h40;
    wire [7:0] \AES.a8_rcon  = 8'h80;
    wire [7:0] \AES.a9_rcon  = 8'h1b;
    wire [7:0] \AES.a10_rcon  = 8'h36;
    wire \AES.a1.clk ;
    wire [127:0] \AES.a1.in ;
    wire [7:0] \AES.a1.rcon ;
    reg [127:0] \AES.a1.out_1 ;
    wire [127:0] \AES.a1.out_2 ;
    wire [31:0] \AES.a1.k0 ;
    wire [31:0] \AES.a1.k1 ;
    wire [31:0] \AES.a1.k2 ;
    wire [31:0] \AES.a1.k3 ;
    wire [31:0] \AES.a1.v0 ;
    wire [31:0] \AES.a1.v1 ;
    wire [31:0] \AES.a1.v2 ;
    wire [31:0] \AES.a1.v3 ;
    reg [31:0] \AES.a1.k0a ;
    reg [31:0] \AES.a1.k1a ;
    reg [31:0] \AES.a1.k2a ;
    reg [31:0] \AES.a1.k3a ;
    wire [31:0] \AES.a1.k0b ;
    wire [31:0] \AES.a1.k1b ;
    wire [31:0] \AES.a1.k2b ;
    wire [31:0] \AES.a1.k3b ;
    wire [31:0] \AES.a1.k4a ;
    wire \AES.a1.S4_0.clk ;
    wire [31:0] \AES.a1.S4_0.in ;
    wire [31:0] \AES.a1.S4_0.out ;
    wire [7:0] \AES.a1.S4_0.k0 ;
    wire [7:0] \AES.a1.S4_0.k1 ;
    wire [7:0] \AES.a1.S4_0.k2 ;
    wire [7:0] \AES.a1.S4_0.k3 ;
    wire \AES.a1.S4_0.S_0.clk ;
    wire [7:0] \AES.a1.S4_0.S_0.in ;
    reg [7:0] \AES.a1.S4_0.S_0.out ;
    wire \AES.a1.S4_0.S_1.clk ;
    wire [7:0] \AES.a1.S4_0.S_1.in ;
    reg [7:0] \AES.a1.S4_0.S_1.out ;
    wire \AES.a1.S4_0.S_2.clk ;
    wire [7:0] \AES.a1.S4_0.S_2.in ;
    reg [7:0] \AES.a1.S4_0.S_2.out ;
    wire \AES.a1.S4_0.S_3.clk ;
    wire [7:0] \AES.a1.S4_0.S_3.in ;
    reg [7:0] \AES.a1.S4_0.S_3.out ;
    wire \AES.a2.clk ;
    wire [127:0] \AES.a2.in ;
    wire [7:0] \AES.a2.rcon ;
    reg [127:0] \AES.a2.out_1 ;
    wire [127:0] \AES.a2.out_2 ;
    wire [31:0] \AES.a2.k0 ;
    wire [31:0] \AES.a2.k1 ;
    wire [31:0] \AES.a2.k2 ;
    wire [31:0] \AES.a2.k3 ;
    wire [31:0] \AES.a2.v0 ;
    wire [31:0] \AES.a2.v1 ;
    wire [31:0] \AES.a2.v2 ;
    wire [31:0] \AES.a2.v3 ;
    reg [31:0] \AES.a2.k0a ;
    reg [31:0] \AES.a2.k1a ;
    reg [31:0] \AES.a2.k2a ;
    reg [31:0] \AES.a2.k3a ;
    wire [31:0] \AES.a2.k0b ;
    wire [31:0] \AES.a2.k1b ;
    wire [31:0] \AES.a2.k2b ;
    wire [31:0] \AES.a2.k3b ;
    wire [31:0] \AES.a2.k4a ;
    wire \AES.a2.S4_0.clk ;
    wire [31:0] \AES.a2.S4_0.in ;
    wire [31:0] \AES.a2.S4_0.out ;
    wire [7:0] \AES.a2.S4_0.k0 ;
    wire [7:0] \AES.a2.S4_0.k1 ;
    wire [7:0] \AES.a2.S4_0.k2 ;
    wire [7:0] \AES.a2.S4_0.k3 ;
    wire \AES.a2.S4_0.S_0.clk ;
    wire [7:0] \AES.a2.S4_0.S_0.in ;
    reg [7:0] \AES.a2.S4_0.S_0.out ;
    wire \AES.a2.S4_0.S_1.clk ;
    wire [7:0] \AES.a2.S4_0.S_1.in ;
    reg [7:0] \AES.a2.S4_0.S_1.out ;
    wire \AES.a2.S4_0.S_2.clk ;
    wire [7:0] \AES.a2.S4_0.S_2.in ;
    reg [7:0] \AES.a2.S4_0.S_2.out ;
    wire \AES.a2.S4_0.S_3.clk ;
    wire [7:0] \AES.a2.S4_0.S_3.in ;
    reg [7:0] \AES.a2.S4_0.S_3.out ;
    wire \AES.a3.clk ;
    wire [127:0] \AES.a3.in ;
    wire [7:0] \AES.a3.rcon ;
    reg [127:0] \AES.a3.out_1 ;
    wire [127:0] \AES.a3.out_2 ;
    wire [31:0] \AES.a3.k0 ;
    wire [31:0] \AES.a3.k1 ;
    wire [31:0] \AES.a3.k2 ;
    wire [31:0] \AES.a3.k3 ;
    wire [31:0] \AES.a3.v0 ;
    wire [31:0] \AES.a3.v1 ;
    wire [31:0] \AES.a3.v2 ;
    wire [31:0] \AES.a3.v3 ;
    reg [31:0] \AES.a3.k0a ;
    reg [31:0] \AES.a3.k1a ;
    reg [31:0] \AES.a3.k2a ;
    reg [31:0] \AES.a3.k3a ;
    wire [31:0] \AES.a3.k0b ;
    wire [31:0] \AES.a3.k1b ;
    wire [31:0] \AES.a3.k2b ;
    wire [31:0] \AES.a3.k3b ;
    wire [31:0] \AES.a3.k4a ;
    wire \AES.a3.S4_0.clk ;
    wire [31:0] \AES.a3.S4_0.in ;
    wire [31:0] \AES.a3.S4_0.out ;
    wire [7:0] \AES.a3.S4_0.k0 ;
    wire [7:0] \AES.a3.S4_0.k1 ;
    wire [7:0] \AES.a3.S4_0.k2 ;
    wire [7:0] \AES.a3.S4_0.k3 ;
    wire \AES.a3.S4_0.S_0.clk ;
    wire [7:0] \AES.a3.S4_0.S_0.in ;
    reg [7:0] \AES.a3.S4_0.S_0.out ;
    wire \AES.a3.S4_0.S_1.clk ;
    wire [7:0] \AES.a3.S4_0.S_1.in ;
    reg [7:0] \AES.a3.S4_0.S_1.out ;
    wire \AES.a3.S4_0.S_2.clk ;
    wire [7:0] \AES.a3.S4_0.S_2.in ;
    reg [7:0] \AES.a3.S4_0.S_2.out ;
    wire \AES.a3.S4_0.S_3.clk ;
    wire [7:0] \AES.a3.S4_0.S_3.in ;
    reg [7:0] \AES.a3.S4_0.S_3.out ;
    wire \AES.a4.clk ;
    wire [127:0] \AES.a4.in ;
    wire [7:0] \AES.a4.rcon ;
    reg [127:0] \AES.a4.out_1 ;
    wire [127:0] \AES.a4.out_2 ;
    wire [31:0] \AES.a4.k0 ;
    wire [31:0] \AES.a4.k1 ;
    wire [31:0] \AES.a4.k2 ;
    wire [31:0] \AES.a4.k3 ;
    wire [31:0] \AES.a4.v0 ;
    wire [31:0] \AES.a4.v1 ;
    wire [31:0] \AES.a4.v2 ;
    wire [31:0] \AES.a4.v3 ;
    reg [31:0] \AES.a4.k0a ;
    reg [31:0] \AES.a4.k1a ;
    reg [31:0] \AES.a4.k2a ;
    reg [31:0] \AES.a4.k3a ;
    wire [31:0] \AES.a4.k0b ;
    wire [31:0] \AES.a4.k1b ;
    wire [31:0] \AES.a4.k2b ;
    wire [31:0] \AES.a4.k3b ;
    wire [31:0] \AES.a4.k4a ;
    wire \AES.a4.S4_0.clk ;
    wire [31:0] \AES.a4.S4_0.in ;
    wire [31:0] \AES.a4.S4_0.out ;
    wire [7:0] \AES.a4.S4_0.k0 ;
    wire [7:0] \AES.a4.S4_0.k1 ;
    wire [7:0] \AES.a4.S4_0.k2 ;
    wire [7:0] \AES.a4.S4_0.k3 ;
    wire \AES.a4.S4_0.S_0.clk ;
    wire [7:0] \AES.a4.S4_0.S_0.in ;
    reg [7:0] \AES.a4.S4_0.S_0.out ;
    wire \AES.a4.S4_0.S_1.clk ;
    wire [7:0] \AES.a4.S4_0.S_1.in ;
    reg [7:0] \AES.a4.S4_0.S_1.out ;
    wire \AES.a4.S4_0.S_2.clk ;
    wire [7:0] \AES.a4.S4_0.S_2.in ;
    reg [7:0] \AES.a4.S4_0.S_2.out ;
    wire \AES.a4.S4_0.S_3.clk ;
    wire [7:0] \AES.a4.S4_0.S_3.in ;
    reg [7:0] \AES.a4.S4_0.S_3.out ;
    wire \AES.a5.clk ;
    wire [127:0] \AES.a5.in ;
    wire [7:0] \AES.a5.rcon ;
    reg [127:0] \AES.a5.out_1 ;
    wire [127:0] \AES.a5.out_2 ;
    wire [31:0] \AES.a5.k0 ;
    wire [31:0] \AES.a5.k1 ;
    wire [31:0] \AES.a5.k2 ;
    wire [31:0] \AES.a5.k3 ;
    wire [31:0] \AES.a5.v0 ;
    wire [31:0] \AES.a5.v1 ;
    wire [31:0] \AES.a5.v2 ;
    wire [31:0] \AES.a5.v3 ;
    reg [31:0] \AES.a5.k0a ;
    reg [31:0] \AES.a5.k1a ;
    reg [31:0] \AES.a5.k2a ;
    reg [31:0] \AES.a5.k3a ;
    wire [31:0] \AES.a5.k0b ;
    wire [31:0] \AES.a5.k1b ;
    wire [31:0] \AES.a5.k2b ;
    wire [31:0] \AES.a5.k3b ;
    wire [31:0] \AES.a5.k4a ;
    wire \AES.a5.S4_0.clk ;
    wire [31:0] \AES.a5.S4_0.in ;
    wire [31:0] \AES.a5.S4_0.out ;
    wire [7:0] \AES.a5.S4_0.k0 ;
    wire [7:0] \AES.a5.S4_0.k1 ;
    wire [7:0] \AES.a5.S4_0.k2 ;
    wire [7:0] \AES.a5.S4_0.k3 ;
    wire \AES.a5.S4_0.S_0.clk ;
    wire [7:0] \AES.a5.S4_0.S_0.in ;
    reg [7:0] \AES.a5.S4_0.S_0.out ;
    wire \AES.a5.S4_0.S_1.clk ;
    wire [7:0] \AES.a5.S4_0.S_1.in ;
    reg [7:0] \AES.a5.S4_0.S_1.out ;
    wire \AES.a5.S4_0.S_2.clk ;
    wire [7:0] \AES.a5.S4_0.S_2.in ;
    reg [7:0] \AES.a5.S4_0.S_2.out ;
    wire \AES.a5.S4_0.S_3.clk ;
    wire [7:0] \AES.a5.S4_0.S_3.in ;
    reg [7:0] \AES.a5.S4_0.S_3.out ;
    wire \AES.a6.clk ;
    wire [127:0] \AES.a6.in ;
    wire [7:0] \AES.a6.rcon ;
    reg [127:0] \AES.a6.out_1 ;
    wire [127:0] \AES.a6.out_2 ;
    wire [31:0] \AES.a6.k0 ;
    wire [31:0] \AES.a6.k1 ;
    wire [31:0] \AES.a6.k2 ;
    wire [31:0] \AES.a6.k3 ;
    wire [31:0] \AES.a6.v0 ;
    wire [31:0] \AES.a6.v1 ;
    wire [31:0] \AES.a6.v2 ;
    wire [31:0] \AES.a6.v3 ;
    reg [31:0] \AES.a6.k0a ;
    reg [31:0] \AES.a6.k1a ;
    reg [31:0] \AES.a6.k2a ;
    reg [31:0] \AES.a6.k3a ;
    wire [31:0] \AES.a6.k0b ;
    wire [31:0] \AES.a6.k1b ;
    wire [31:0] \AES.a6.k2b ;
    wire [31:0] \AES.a6.k3b ;
    wire [31:0] \AES.a6.k4a ;
    wire \AES.a6.S4_0.clk ;
    wire [31:0] \AES.a6.S4_0.in ;
    wire [31:0] \AES.a6.S4_0.out ;
    wire [7:0] \AES.a6.S4_0.k0 ;
    wire [7:0] \AES.a6.S4_0.k1 ;
    wire [7:0] \AES.a6.S4_0.k2 ;
    wire [7:0] \AES.a6.S4_0.k3 ;
    wire \AES.a6.S4_0.S_0.clk ;
    wire [7:0] \AES.a6.S4_0.S_0.in ;
    reg [7:0] \AES.a6.S4_0.S_0.out ;
    wire \AES.a6.S4_0.S_1.clk ;
    wire [7:0] \AES.a6.S4_0.S_1.in ;
    reg [7:0] \AES.a6.S4_0.S_1.out ;
    wire \AES.a6.S4_0.S_2.clk ;
    wire [7:0] \AES.a6.S4_0.S_2.in ;
    reg [7:0] \AES.a6.S4_0.S_2.out ;
    wire \AES.a6.S4_0.S_3.clk ;
    wire [7:0] \AES.a6.S4_0.S_3.in ;
    reg [7:0] \AES.a6.S4_0.S_3.out ;
    wire \AES.a7.clk ;
    wire [127:0] \AES.a7.in ;
    wire [7:0] \AES.a7.rcon ;
    reg [127:0] \AES.a7.out_1 ;
    wire [127:0] \AES.a7.out_2 ;
    wire [31:0] \AES.a7.k0 ;
    wire [31:0] \AES.a7.k1 ;
    wire [31:0] \AES.a7.k2 ;
    wire [31:0] \AES.a7.k3 ;
    wire [31:0] \AES.a7.v0 ;
    wire [31:0] \AES.a7.v1 ;
    wire [31:0] \AES.a7.v2 ;
    wire [31:0] \AES.a7.v3 ;
    reg [31:0] \AES.a7.k0a ;
    reg [31:0] \AES.a7.k1a ;
    reg [31:0] \AES.a7.k2a ;
    reg [31:0] \AES.a7.k3a ;
    wire [31:0] \AES.a7.k0b ;
    wire [31:0] \AES.a7.k1b ;
    wire [31:0] \AES.a7.k2b ;
    wire [31:0] \AES.a7.k3b ;
    wire [31:0] \AES.a7.k4a ;
    wire \AES.a7.S4_0.clk ;
    wire [31:0] \AES.a7.S4_0.in ;
    wire [31:0] \AES.a7.S4_0.out ;
    wire [7:0] \AES.a7.S4_0.k0 ;
    wire [7:0] \AES.a7.S4_0.k1 ;
    wire [7:0] \AES.a7.S4_0.k2 ;
    wire [7:0] \AES.a7.S4_0.k3 ;
    wire \AES.a7.S4_0.S_0.clk ;
    wire [7:0] \AES.a7.S4_0.S_0.in ;
    reg [7:0] \AES.a7.S4_0.S_0.out ;
    wire \AES.a7.S4_0.S_1.clk ;
    wire [7:0] \AES.a7.S4_0.S_1.in ;
    reg [7:0] \AES.a7.S4_0.S_1.out ;
    wire \AES.a7.S4_0.S_2.clk ;
    wire [7:0] \AES.a7.S4_0.S_2.in ;
    reg [7:0] \AES.a7.S4_0.S_2.out ;
    wire \AES.a7.S4_0.S_3.clk ;
    wire [7:0] \AES.a7.S4_0.S_3.in ;
    reg [7:0] \AES.a7.S4_0.S_3.out ;
    wire \AES.a8.clk ;
    wire [127:0] \AES.a8.in ;
    wire [7:0] \AES.a8.rcon ;
    reg [127:0] \AES.a8.out_1 ;
    wire [127:0] \AES.a8.out_2 ;
    wire [31:0] \AES.a8.k0 ;
    wire [31:0] \AES.a8.k1 ;
    wire [31:0] \AES.a8.k2 ;
    wire [31:0] \AES.a8.k3 ;
    wire [31:0] \AES.a8.v0 ;
    wire [31:0] \AES.a8.v1 ;
    wire [31:0] \AES.a8.v2 ;
    wire [31:0] \AES.a8.v3 ;
    reg [31:0] \AES.a8.k0a ;
    reg [31:0] \AES.a8.k1a ;
    reg [31:0] \AES.a8.k2a ;
    reg [31:0] \AES.a8.k3a ;
    wire [31:0] \AES.a8.k0b ;
    wire [31:0] \AES.a8.k1b ;
    wire [31:0] \AES.a8.k2b ;
    wire [31:0] \AES.a8.k3b ;
    wire [31:0] \AES.a8.k4a ;
    wire \AES.a8.S4_0.clk ;
    wire [31:0] \AES.a8.S4_0.in ;
    wire [31:0] \AES.a8.S4_0.out ;
    wire [7:0] \AES.a8.S4_0.k0 ;
    wire [7:0] \AES.a8.S4_0.k1 ;
    wire [7:0] \AES.a8.S4_0.k2 ;
    wire [7:0] \AES.a8.S4_0.k3 ;
    wire \AES.a8.S4_0.S_0.clk ;
    wire [7:0] \AES.a8.S4_0.S_0.in ;
    reg [7:0] \AES.a8.S4_0.S_0.out ;
    wire \AES.a8.S4_0.S_1.clk ;
    wire [7:0] \AES.a8.S4_0.S_1.in ;
    reg [7:0] \AES.a8.S4_0.S_1.out ;
    wire \AES.a8.S4_0.S_2.clk ;
    wire [7:0] \AES.a8.S4_0.S_2.in ;
    reg [7:0] \AES.a8.S4_0.S_2.out ;
    wire \AES.a8.S4_0.S_3.clk ;
    wire [7:0] \AES.a8.S4_0.S_3.in ;
    reg [7:0] \AES.a8.S4_0.S_3.out ;
    wire \AES.a9.clk ;
    wire [127:0] \AES.a9.in ;
    wire [7:0] \AES.a9.rcon ;
    reg [127:0] \AES.a9.out_1 ;
    wire [127:0] \AES.a9.out_2 ;
    wire [31:0] \AES.a9.k0 ;
    wire [31:0] \AES.a9.k1 ;
    wire [31:0] \AES.a9.k2 ;
    wire [31:0] \AES.a9.k3 ;
    wire [31:0] \AES.a9.v0 ;
    wire [31:0] \AES.a9.v1 ;
    wire [31:0] \AES.a9.v2 ;
    wire [31:0] \AES.a9.v3 ;
    reg [31:0] \AES.a9.k0a ;
    reg [31:0] \AES.a9.k1a ;
    reg [31:0] \AES.a9.k2a ;
    reg [31:0] \AES.a9.k3a ;
    wire [31:0] \AES.a9.k0b ;
    wire [31:0] \AES.a9.k1b ;
    wire [31:0] \AES.a9.k2b ;
    wire [31:0] \AES.a9.k3b ;
    wire [31:0] \AES.a9.k4a ;
    wire \AES.a9.S4_0.clk ;
    wire [31:0] \AES.a9.S4_0.in ;
    wire [31:0] \AES.a9.S4_0.out ;
    wire [7:0] \AES.a9.S4_0.k0 ;
    wire [7:0] \AES.a9.S4_0.k1 ;
    wire [7:0] \AES.a9.S4_0.k2 ;
    wire [7:0] \AES.a9.S4_0.k3 ;
    wire \AES.a9.S4_0.S_0.clk ;
    wire [7:0] \AES.a9.S4_0.S_0.in ;
    reg [7:0] \AES.a9.S4_0.S_0.out ;
    wire \AES.a9.S4_0.S_1.clk ;
    wire [7:0] \AES.a9.S4_0.S_1.in ;
    reg [7:0] \AES.a9.S4_0.S_1.out ;
    wire \AES.a9.S4_0.S_2.clk ;
    wire [7:0] \AES.a9.S4_0.S_2.in ;
    reg [7:0] \AES.a9.S4_0.S_2.out ;
    wire \AES.a9.S4_0.S_3.clk ;
    wire [7:0] \AES.a9.S4_0.S_3.in ;
    reg [7:0] \AES.a9.S4_0.S_3.out ;
    wire \AES.a10.clk ;
    wire [127:0] \AES.a10.in ;
    wire [7:0] \AES.a10.rcon ;
    reg [127:0] \AES.a10.out_1 ;
    wire [127:0] \AES.a10.out_2 ;
    wire [31:0] \AES.a10.k0 ;
    wire [31:0] \AES.a10.k1 ;
    wire [31:0] \AES.a10.k2 ;
    wire [31:0] \AES.a10.k3 ;
    wire [31:0] \AES.a10.v0 ;
    wire [31:0] \AES.a10.v1 ;
    wire [31:0] \AES.a10.v2 ;
    wire [31:0] \AES.a10.v3 ;
    reg [31:0] \AES.a10.k0a ;
    reg [31:0] \AES.a10.k1a ;
    reg [31:0] \AES.a10.k2a ;
    reg [31:0] \AES.a10.k3a ;
    wire [31:0] \AES.a10.k0b ;
    wire [31:0] \AES.a10.k1b ;
    wire [31:0] \AES.a10.k2b ;
    wire [31:0] \AES.a10.k3b ;
    wire [31:0] \AES.a10.k4a ;
    wire \AES.a10.S4_0.clk ;
    wire [31:0] \AES.a10.S4_0.in ;
    wire [31:0] \AES.a10.S4_0.out ;
    wire [7:0] \AES.a10.S4_0.k0 ;
    wire [7:0] \AES.a10.S4_0.k1 ;
    wire [7:0] \AES.a10.S4_0.k2 ;
    wire [7:0] \AES.a10.S4_0.k3 ;
    wire \AES.a10.S4_0.S_0.clk ;
    wire [7:0] \AES.a10.S4_0.S_0.in ;
    reg [7:0] \AES.a10.S4_0.S_0.out ;
    wire \AES.a10.S4_0.S_1.clk ;
    wire [7:0] \AES.a10.S4_0.S_1.in ;
    reg [7:0] \AES.a10.S4_0.S_1.out ;
    wire \AES.a10.S4_0.S_2.clk ;
    wire [7:0] \AES.a10.S4_0.S_2.in ;
    reg [7:0] \AES.a10.S4_0.S_2.out ;
    wire \AES.a10.S4_0.S_3.clk ;
    wire [7:0] \AES.a10.S4_0.S_3.in ;
    reg [7:0] \AES.a10.S4_0.S_3.out ;
    wire \AES.r1.clk ;
    wire [127:0] \AES.r1.state_in ;
    wire [127:0] \AES.r1.key ;
    reg [127:0] \AES.r1.state_out ;
    wire [31:0] \AES.r1.s0 ;
    wire [31:0] \AES.r1.s1 ;
    wire [31:0] \AES.r1.s2 ;
    wire [31:0] \AES.r1.s3 ;
    wire [31:0] \AES.r1.z0 ;
    wire [31:0] \AES.r1.z1 ;
    wire [31:0] \AES.r1.z2 ;
    wire [31:0] \AES.r1.z3 ;
    wire [31:0] \AES.r1.p00 ;
    wire [31:0] \AES.r1.p01 ;
    wire [31:0] \AES.r1.p02 ;
    wire [31:0] \AES.r1.p03 ;
    wire [31:0] \AES.r1.p10 ;
    wire [31:0] \AES.r1.p11 ;
    wire [31:0] \AES.r1.p12 ;
    wire [31:0] \AES.r1.p13 ;
    wire [31:0] \AES.r1.p20 ;
    wire [31:0] \AES.r1.p21 ;
    wire [31:0] \AES.r1.p22 ;
    wire [31:0] \AES.r1.p23 ;
    wire [31:0] \AES.r1.p30 ;
    wire [31:0] \AES.r1.p31 ;
    wire [31:0] \AES.r1.p32 ;
    wire [31:0] \AES.r1.p33 ;
    wire [31:0] \AES.r1.k0 ;
    wire [31:0] \AES.r1.k1 ;
    wire [31:0] \AES.r1.k2 ;
    wire [31:0] \AES.r1.k3 ;
    wire \AES.r1.t0.clk ;
    wire [31:0] \AES.r1.t0.state ;
    wire [31:0] \AES.r1.t0.p0 ;
    wire [31:0] \AES.r1.t0.p1 ;
    wire [31:0] \AES.r1.t0.p2 ;
    wire [31:0] \AES.r1.t0.p3 ;
    wire [7:0] \AES.r1.t0.b0 ;
    wire [7:0] \AES.r1.t0.b1 ;
    wire [7:0] \AES.r1.t0.b2 ;
    wire [7:0] \AES.r1.t0.b3 ;
    wire [31:0] \AES.r1.t0.k0 ;
    wire [31:0] \AES.r1.t0.k1 ;
    wire [31:0] \AES.r1.t0.k2 ;
    wire \AES.r1.t0.t0.clk ;
    wire [7:0] \AES.r1.t0.t0.in ;
    wire [31:0] \AES.r1.t0.t0.out ;
    wire [7:0] \AES.r1.t0.t0.k0 ;
    wire [7:0] \AES.r1.t0.t0.k1 ;
    wire \AES.r1.t0.t0.s0.clk ;
    wire [7:0] \AES.r1.t0.t0.s0.in ;
    reg [7:0] \AES.r1.t0.t0.s0.out ;
    wire \AES.r1.t0.t0.s4.clk ;
    wire [7:0] \AES.r1.t0.t0.s4.in ;
    reg [7:0] \AES.r1.t0.t0.s4.out ;
    wire \AES.r1.t0.t1.clk ;
    wire [7:0] \AES.r1.t0.t1.in ;
    wire [31:0] \AES.r1.t0.t1.out ;
    wire [7:0] \AES.r1.t0.t1.k0 ;
    wire [7:0] \AES.r1.t0.t1.k1 ;
    wire \AES.r1.t0.t1.s0.clk ;
    wire [7:0] \AES.r1.t0.t1.s0.in ;
    reg [7:0] \AES.r1.t0.t1.s0.out ;
    wire \AES.r1.t0.t1.s4.clk ;
    wire [7:0] \AES.r1.t0.t1.s4.in ;
    reg [7:0] \AES.r1.t0.t1.s4.out ;
    wire \AES.r1.t0.t2.clk ;
    wire [7:0] \AES.r1.t0.t2.in ;
    wire [31:0] \AES.r1.t0.t2.out ;
    wire [7:0] \AES.r1.t0.t2.k0 ;
    wire [7:0] \AES.r1.t0.t2.k1 ;
    wire \AES.r1.t0.t2.s0.clk ;
    wire [7:0] \AES.r1.t0.t2.s0.in ;
    reg [7:0] \AES.r1.t0.t2.s0.out ;
    wire \AES.r1.t0.t2.s4.clk ;
    wire [7:0] \AES.r1.t0.t2.s4.in ;
    reg [7:0] \AES.r1.t0.t2.s4.out ;
    wire \AES.r1.t0.t3.clk ;
    wire [7:0] \AES.r1.t0.t3.in ;
    wire [31:0] \AES.r1.t0.t3.out ;
    wire [7:0] \AES.r1.t0.t3.k0 ;
    wire [7:0] \AES.r1.t0.t3.k1 ;
    wire \AES.r1.t0.t3.s0.clk ;
    wire [7:0] \AES.r1.t0.t3.s0.in ;
    reg [7:0] \AES.r1.t0.t3.s0.out ;
    wire \AES.r1.t0.t3.s4.clk ;
    wire [7:0] \AES.r1.t0.t3.s4.in ;
    reg [7:0] \AES.r1.t0.t3.s4.out ;
    wire \AES.r1.t1.clk ;
    wire [31:0] \AES.r1.t1.state ;
    wire [31:0] \AES.r1.t1.p0 ;
    wire [31:0] \AES.r1.t1.p1 ;
    wire [31:0] \AES.r1.t1.p2 ;
    wire [31:0] \AES.r1.t1.p3 ;
    wire [7:0] \AES.r1.t1.b0 ;
    wire [7:0] \AES.r1.t1.b1 ;
    wire [7:0] \AES.r1.t1.b2 ;
    wire [7:0] \AES.r1.t1.b3 ;
    wire [31:0] \AES.r1.t1.k0 ;
    wire [31:0] \AES.r1.t1.k1 ;
    wire [31:0] \AES.r1.t1.k2 ;
    wire \AES.r1.t1.t0.clk ;
    wire [7:0] \AES.r1.t1.t0.in ;
    wire [31:0] \AES.r1.t1.t0.out ;
    wire [7:0] \AES.r1.t1.t0.k0 ;
    wire [7:0] \AES.r1.t1.t0.k1 ;
    wire \AES.r1.t1.t0.s0.clk ;
    wire [7:0] \AES.r1.t1.t0.s0.in ;
    reg [7:0] \AES.r1.t1.t0.s0.out ;
    wire \AES.r1.t1.t0.s4.clk ;
    wire [7:0] \AES.r1.t1.t0.s4.in ;
    reg [7:0] \AES.r1.t1.t0.s4.out ;
    wire \AES.r1.t1.t1.clk ;
    wire [7:0] \AES.r1.t1.t1.in ;
    wire [31:0] \AES.r1.t1.t1.out ;
    wire [7:0] \AES.r1.t1.t1.k0 ;
    wire [7:0] \AES.r1.t1.t1.k1 ;
    wire \AES.r1.t1.t1.s0.clk ;
    wire [7:0] \AES.r1.t1.t1.s0.in ;
    reg [7:0] \AES.r1.t1.t1.s0.out ;
    wire \AES.r1.t1.t1.s4.clk ;
    wire [7:0] \AES.r1.t1.t1.s4.in ;
    reg [7:0] \AES.r1.t1.t1.s4.out ;
    wire \AES.r1.t1.t2.clk ;
    wire [7:0] \AES.r1.t1.t2.in ;
    wire [31:0] \AES.r1.t1.t2.out ;
    wire [7:0] \AES.r1.t1.t2.k0 ;
    wire [7:0] \AES.r1.t1.t2.k1 ;
    wire \AES.r1.t1.t2.s0.clk ;
    wire [7:0] \AES.r1.t1.t2.s0.in ;
    reg [7:0] \AES.r1.t1.t2.s0.out ;
    wire \AES.r1.t1.t2.s4.clk ;
    wire [7:0] \AES.r1.t1.t2.s4.in ;
    reg [7:0] \AES.r1.t1.t2.s4.out ;
    wire \AES.r1.t1.t3.clk ;
    wire [7:0] \AES.r1.t1.t3.in ;
    wire [31:0] \AES.r1.t1.t3.out ;
    wire [7:0] \AES.r1.t1.t3.k0 ;
    wire [7:0] \AES.r1.t1.t3.k1 ;
    wire \AES.r1.t1.t3.s0.clk ;
    wire [7:0] \AES.r1.t1.t3.s0.in ;
    reg [7:0] \AES.r1.t1.t3.s0.out ;
    wire \AES.r1.t1.t3.s4.clk ;
    wire [7:0] \AES.r1.t1.t3.s4.in ;
    reg [7:0] \AES.r1.t1.t3.s4.out ;
    wire \AES.r1.t2.clk ;
    wire [31:0] \AES.r1.t2.state ;
    wire [31:0] \AES.r1.t2.p0 ;
    wire [31:0] \AES.r1.t2.p1 ;
    wire [31:0] \AES.r1.t2.p2 ;
    wire [31:0] \AES.r1.t2.p3 ;
    wire [7:0] \AES.r1.t2.b0 ;
    wire [7:0] \AES.r1.t2.b1 ;
    wire [7:0] \AES.r1.t2.b2 ;
    wire [7:0] \AES.r1.t2.b3 ;
    wire [31:0] \AES.r1.t2.k0 ;
    wire [31:0] \AES.r1.t2.k1 ;
    wire [31:0] \AES.r1.t2.k2 ;
    wire \AES.r1.t2.t0.clk ;
    wire [7:0] \AES.r1.t2.t0.in ;
    wire [31:0] \AES.r1.t2.t0.out ;
    wire [7:0] \AES.r1.t2.t0.k0 ;
    wire [7:0] \AES.r1.t2.t0.k1 ;
    wire \AES.r1.t2.t0.s0.clk ;
    wire [7:0] \AES.r1.t2.t0.s0.in ;
    reg [7:0] \AES.r1.t2.t0.s0.out ;
    wire \AES.r1.t2.t0.s4.clk ;
    wire [7:0] \AES.r1.t2.t0.s4.in ;
    reg [7:0] \AES.r1.t2.t0.s4.out ;
    wire \AES.r1.t2.t1.clk ;
    wire [7:0] \AES.r1.t2.t1.in ;
    wire [31:0] \AES.r1.t2.t1.out ;
    wire [7:0] \AES.r1.t2.t1.k0 ;
    wire [7:0] \AES.r1.t2.t1.k1 ;
    wire \AES.r1.t2.t1.s0.clk ;
    wire [7:0] \AES.r1.t2.t1.s0.in ;
    reg [7:0] \AES.r1.t2.t1.s0.out ;
    wire \AES.r1.t2.t1.s4.clk ;
    wire [7:0] \AES.r1.t2.t1.s4.in ;
    reg [7:0] \AES.r1.t2.t1.s4.out ;
    wire \AES.r1.t2.t2.clk ;
    wire [7:0] \AES.r1.t2.t2.in ;
    wire [31:0] \AES.r1.t2.t2.out ;
    wire [7:0] \AES.r1.t2.t2.k0 ;
    wire [7:0] \AES.r1.t2.t2.k1 ;
    wire \AES.r1.t2.t2.s0.clk ;
    wire [7:0] \AES.r1.t2.t2.s0.in ;
    reg [7:0] \AES.r1.t2.t2.s0.out ;
    wire \AES.r1.t2.t2.s4.clk ;
    wire [7:0] \AES.r1.t2.t2.s4.in ;
    reg [7:0] \AES.r1.t2.t2.s4.out ;
    wire \AES.r1.t2.t3.clk ;
    wire [7:0] \AES.r1.t2.t3.in ;
    wire [31:0] \AES.r1.t2.t3.out ;
    wire [7:0] \AES.r1.t2.t3.k0 ;
    wire [7:0] \AES.r1.t2.t3.k1 ;
    wire \AES.r1.t2.t3.s0.clk ;
    wire [7:0] \AES.r1.t2.t3.s0.in ;
    reg [7:0] \AES.r1.t2.t3.s0.out ;
    wire \AES.r1.t2.t3.s4.clk ;
    wire [7:0] \AES.r1.t2.t3.s4.in ;
    reg [7:0] \AES.r1.t2.t3.s4.out ;
    wire \AES.r1.t3.clk ;
    wire [31:0] \AES.r1.t3.state ;
    wire [31:0] \AES.r1.t3.p0 ;
    wire [31:0] \AES.r1.t3.p1 ;
    wire [31:0] \AES.r1.t3.p2 ;
    wire [31:0] \AES.r1.t3.p3 ;
    wire [7:0] \AES.r1.t3.b0 ;
    wire [7:0] \AES.r1.t3.b1 ;
    wire [7:0] \AES.r1.t3.b2 ;
    wire [7:0] \AES.r1.t3.b3 ;
    wire [31:0] \AES.r1.t3.k0 ;
    wire [31:0] \AES.r1.t3.k1 ;
    wire [31:0] \AES.r1.t3.k2 ;
    wire \AES.r1.t3.t0.clk ;
    wire [7:0] \AES.r1.t3.t0.in ;
    wire [31:0] \AES.r1.t3.t0.out ;
    wire [7:0] \AES.r1.t3.t0.k0 ;
    wire [7:0] \AES.r1.t3.t0.k1 ;
    wire \AES.r1.t3.t0.s0.clk ;
    wire [7:0] \AES.r1.t3.t0.s0.in ;
    reg [7:0] \AES.r1.t3.t0.s0.out ;
    wire \AES.r1.t3.t0.s4.clk ;
    wire [7:0] \AES.r1.t3.t0.s4.in ;
    reg [7:0] \AES.r1.t3.t0.s4.out ;
    wire \AES.r1.t3.t1.clk ;
    wire [7:0] \AES.r1.t3.t1.in ;
    wire [31:0] \AES.r1.t3.t1.out ;
    wire [7:0] \AES.r1.t3.t1.k0 ;
    wire [7:0] \AES.r1.t3.t1.k1 ;
    wire \AES.r1.t3.t1.s0.clk ;
    wire [7:0] \AES.r1.t3.t1.s0.in ;
    reg [7:0] \AES.r1.t3.t1.s0.out ;
    wire \AES.r1.t3.t1.s4.clk ;
    wire [7:0] \AES.r1.t3.t1.s4.in ;
    reg [7:0] \AES.r1.t3.t1.s4.out ;
    wire \AES.r1.t3.t2.clk ;
    wire [7:0] \AES.r1.t3.t2.in ;
    wire [31:0] \AES.r1.t3.t2.out ;
    wire [7:0] \AES.r1.t3.t2.k0 ;
    wire [7:0] \AES.r1.t3.t2.k1 ;
    wire \AES.r1.t3.t2.s0.clk ;
    wire [7:0] \AES.r1.t3.t2.s0.in ;
    reg [7:0] \AES.r1.t3.t2.s0.out ;
    wire \AES.r1.t3.t2.s4.clk ;
    wire [7:0] \AES.r1.t3.t2.s4.in ;
    reg [7:0] \AES.r1.t3.t2.s4.out ;
    wire \AES.r1.t3.t3.clk ;
    wire [7:0] \AES.r1.t3.t3.in ;
    wire [31:0] \AES.r1.t3.t3.out ;
    wire [7:0] \AES.r1.t3.t3.k0 ;
    wire [7:0] \AES.r1.t3.t3.k1 ;
    wire \AES.r1.t3.t3.s0.clk ;
    wire [7:0] \AES.r1.t3.t3.s0.in ;
    reg [7:0] \AES.r1.t3.t3.s0.out ;
    wire \AES.r1.t3.t3.s4.clk ;
    wire [7:0] \AES.r1.t3.t3.s4.in ;
    reg [7:0] \AES.r1.t3.t3.s4.out ;
    wire \AES.r2.clk ;
    wire [127:0] \AES.r2.state_in ;
    wire [127:0] \AES.r2.key ;
    reg [127:0] \AES.r2.state_out ;
    wire [31:0] \AES.r2.s0 ;
    wire [31:0] \AES.r2.s1 ;
    wire [31:0] \AES.r2.s2 ;
    wire [31:0] \AES.r2.s3 ;
    wire [31:0] \AES.r2.z0 ;
    wire [31:0] \AES.r2.z1 ;
    wire [31:0] \AES.r2.z2 ;
    wire [31:0] \AES.r2.z3 ;
    wire [31:0] \AES.r2.p00 ;
    wire [31:0] \AES.r2.p01 ;
    wire [31:0] \AES.r2.p02 ;
    wire [31:0] \AES.r2.p03 ;
    wire [31:0] \AES.r2.p10 ;
    wire [31:0] \AES.r2.p11 ;
    wire [31:0] \AES.r2.p12 ;
    wire [31:0] \AES.r2.p13 ;
    wire [31:0] \AES.r2.p20 ;
    wire [31:0] \AES.r2.p21 ;
    wire [31:0] \AES.r2.p22 ;
    wire [31:0] \AES.r2.p23 ;
    wire [31:0] \AES.r2.p30 ;
    wire [31:0] \AES.r2.p31 ;
    wire [31:0] \AES.r2.p32 ;
    wire [31:0] \AES.r2.p33 ;
    wire [31:0] \AES.r2.k0 ;
    wire [31:0] \AES.r2.k1 ;
    wire [31:0] \AES.r2.k2 ;
    wire [31:0] \AES.r2.k3 ;
    wire \AES.r2.t0.clk ;
    wire [31:0] \AES.r2.t0.state ;
    wire [31:0] \AES.r2.t0.p0 ;
    wire [31:0] \AES.r2.t0.p1 ;
    wire [31:0] \AES.r2.t0.p2 ;
    wire [31:0] \AES.r2.t0.p3 ;
    wire [7:0] \AES.r2.t0.b0 ;
    wire [7:0] \AES.r2.t0.b1 ;
    wire [7:0] \AES.r2.t0.b2 ;
    wire [7:0] \AES.r2.t0.b3 ;
    wire [31:0] \AES.r2.t0.k0 ;
    wire [31:0] \AES.r2.t0.k1 ;
    wire [31:0] \AES.r2.t0.k2 ;
    wire \AES.r2.t0.t0.clk ;
    wire [7:0] \AES.r2.t0.t0.in ;
    wire [31:0] \AES.r2.t0.t0.out ;
    wire [7:0] \AES.r2.t0.t0.k0 ;
    wire [7:0] \AES.r2.t0.t0.k1 ;
    wire \AES.r2.t0.t0.s0.clk ;
    wire [7:0] \AES.r2.t0.t0.s0.in ;
    reg [7:0] \AES.r2.t0.t0.s0.out ;
    wire \AES.r2.t0.t0.s4.clk ;
    wire [7:0] \AES.r2.t0.t0.s4.in ;
    reg [7:0] \AES.r2.t0.t0.s4.out ;
    wire \AES.r2.t0.t1.clk ;
    wire [7:0] \AES.r2.t0.t1.in ;
    wire [31:0] \AES.r2.t0.t1.out ;
    wire [7:0] \AES.r2.t0.t1.k0 ;
    wire [7:0] \AES.r2.t0.t1.k1 ;
    wire \AES.r2.t0.t1.s0.clk ;
    wire [7:0] \AES.r2.t0.t1.s0.in ;
    reg [7:0] \AES.r2.t0.t1.s0.out ;
    wire \AES.r2.t0.t1.s4.clk ;
    wire [7:0] \AES.r2.t0.t1.s4.in ;
    reg [7:0] \AES.r2.t0.t1.s4.out ;
    wire \AES.r2.t0.t2.clk ;
    wire [7:0] \AES.r2.t0.t2.in ;
    wire [31:0] \AES.r2.t0.t2.out ;
    wire [7:0] \AES.r2.t0.t2.k0 ;
    wire [7:0] \AES.r2.t0.t2.k1 ;
    wire \AES.r2.t0.t2.s0.clk ;
    wire [7:0] \AES.r2.t0.t2.s0.in ;
    reg [7:0] \AES.r2.t0.t2.s0.out ;
    wire \AES.r2.t0.t2.s4.clk ;
    wire [7:0] \AES.r2.t0.t2.s4.in ;
    reg [7:0] \AES.r2.t0.t2.s4.out ;
    wire \AES.r2.t0.t3.clk ;
    wire [7:0] \AES.r2.t0.t3.in ;
    wire [31:0] \AES.r2.t0.t3.out ;
    wire [7:0] \AES.r2.t0.t3.k0 ;
    wire [7:0] \AES.r2.t0.t3.k1 ;
    wire \AES.r2.t0.t3.s0.clk ;
    wire [7:0] \AES.r2.t0.t3.s0.in ;
    reg [7:0] \AES.r2.t0.t3.s0.out ;
    wire \AES.r2.t0.t3.s4.clk ;
    wire [7:0] \AES.r2.t0.t3.s4.in ;
    reg [7:0] \AES.r2.t0.t3.s4.out ;
    wire \AES.r2.t1.clk ;
    wire [31:0] \AES.r2.t1.state ;
    wire [31:0] \AES.r2.t1.p0 ;
    wire [31:0] \AES.r2.t1.p1 ;
    wire [31:0] \AES.r2.t1.p2 ;
    wire [31:0] \AES.r2.t1.p3 ;
    wire [7:0] \AES.r2.t1.b0 ;
    wire [7:0] \AES.r2.t1.b1 ;
    wire [7:0] \AES.r2.t1.b2 ;
    wire [7:0] \AES.r2.t1.b3 ;
    wire [31:0] \AES.r2.t1.k0 ;
    wire [31:0] \AES.r2.t1.k1 ;
    wire [31:0] \AES.r2.t1.k2 ;
    wire \AES.r2.t1.t0.clk ;
    wire [7:0] \AES.r2.t1.t0.in ;
    wire [31:0] \AES.r2.t1.t0.out ;
    wire [7:0] \AES.r2.t1.t0.k0 ;
    wire [7:0] \AES.r2.t1.t0.k1 ;
    wire \AES.r2.t1.t0.s0.clk ;
    wire [7:0] \AES.r2.t1.t0.s0.in ;
    reg [7:0] \AES.r2.t1.t0.s0.out ;
    wire \AES.r2.t1.t0.s4.clk ;
    wire [7:0] \AES.r2.t1.t0.s4.in ;
    reg [7:0] \AES.r2.t1.t0.s4.out ;
    wire \AES.r2.t1.t1.clk ;
    wire [7:0] \AES.r2.t1.t1.in ;
    wire [31:0] \AES.r2.t1.t1.out ;
    wire [7:0] \AES.r2.t1.t1.k0 ;
    wire [7:0] \AES.r2.t1.t1.k1 ;
    wire \AES.r2.t1.t1.s0.clk ;
    wire [7:0] \AES.r2.t1.t1.s0.in ;
    reg [7:0] \AES.r2.t1.t1.s0.out ;
    wire \AES.r2.t1.t1.s4.clk ;
    wire [7:0] \AES.r2.t1.t1.s4.in ;
    reg [7:0] \AES.r2.t1.t1.s4.out ;
    wire \AES.r2.t1.t2.clk ;
    wire [7:0] \AES.r2.t1.t2.in ;
    wire [31:0] \AES.r2.t1.t2.out ;
    wire [7:0] \AES.r2.t1.t2.k0 ;
    wire [7:0] \AES.r2.t1.t2.k1 ;
    wire \AES.r2.t1.t2.s0.clk ;
    wire [7:0] \AES.r2.t1.t2.s0.in ;
    reg [7:0] \AES.r2.t1.t2.s0.out ;
    wire \AES.r2.t1.t2.s4.clk ;
    wire [7:0] \AES.r2.t1.t2.s4.in ;
    reg [7:0] \AES.r2.t1.t2.s4.out ;
    wire \AES.r2.t1.t3.clk ;
    wire [7:0] \AES.r2.t1.t3.in ;
    wire [31:0] \AES.r2.t1.t3.out ;
    wire [7:0] \AES.r2.t1.t3.k0 ;
    wire [7:0] \AES.r2.t1.t3.k1 ;
    wire \AES.r2.t1.t3.s0.clk ;
    wire [7:0] \AES.r2.t1.t3.s0.in ;
    reg [7:0] \AES.r2.t1.t3.s0.out ;
    wire \AES.r2.t1.t3.s4.clk ;
    wire [7:0] \AES.r2.t1.t3.s4.in ;
    reg [7:0] \AES.r2.t1.t3.s4.out ;
    wire \AES.r2.t2.clk ;
    wire [31:0] \AES.r2.t2.state ;
    wire [31:0] \AES.r2.t2.p0 ;
    wire [31:0] \AES.r2.t2.p1 ;
    wire [31:0] \AES.r2.t2.p2 ;
    wire [31:0] \AES.r2.t2.p3 ;
    wire [7:0] \AES.r2.t2.b0 ;
    wire [7:0] \AES.r2.t2.b1 ;
    wire [7:0] \AES.r2.t2.b2 ;
    wire [7:0] \AES.r2.t2.b3 ;
    wire [31:0] \AES.r2.t2.k0 ;
    wire [31:0] \AES.r2.t2.k1 ;
    wire [31:0] \AES.r2.t2.k2 ;
    wire \AES.r2.t2.t0.clk ;
    wire [7:0] \AES.r2.t2.t0.in ;
    wire [31:0] \AES.r2.t2.t0.out ;
    wire [7:0] \AES.r2.t2.t0.k0 ;
    wire [7:0] \AES.r2.t2.t0.k1 ;
    wire \AES.r2.t2.t0.s0.clk ;
    wire [7:0] \AES.r2.t2.t0.s0.in ;
    reg [7:0] \AES.r2.t2.t0.s0.out ;
    wire \AES.r2.t2.t0.s4.clk ;
    wire [7:0] \AES.r2.t2.t0.s4.in ;
    reg [7:0] \AES.r2.t2.t0.s4.out ;
    wire \AES.r2.t2.t1.clk ;
    wire [7:0] \AES.r2.t2.t1.in ;
    wire [31:0] \AES.r2.t2.t1.out ;
    wire [7:0] \AES.r2.t2.t1.k0 ;
    wire [7:0] \AES.r2.t2.t1.k1 ;
    wire \AES.r2.t2.t1.s0.clk ;
    wire [7:0] \AES.r2.t2.t1.s0.in ;
    reg [7:0] \AES.r2.t2.t1.s0.out ;
    wire \AES.r2.t2.t1.s4.clk ;
    wire [7:0] \AES.r2.t2.t1.s4.in ;
    reg [7:0] \AES.r2.t2.t1.s4.out ;
    wire \AES.r2.t2.t2.clk ;
    wire [7:0] \AES.r2.t2.t2.in ;
    wire [31:0] \AES.r2.t2.t2.out ;
    wire [7:0] \AES.r2.t2.t2.k0 ;
    wire [7:0] \AES.r2.t2.t2.k1 ;
    wire \AES.r2.t2.t2.s0.clk ;
    wire [7:0] \AES.r2.t2.t2.s0.in ;
    reg [7:0] \AES.r2.t2.t2.s0.out ;
    wire \AES.r2.t2.t2.s4.clk ;
    wire [7:0] \AES.r2.t2.t2.s4.in ;
    reg [7:0] \AES.r2.t2.t2.s4.out ;
    wire \AES.r2.t2.t3.clk ;
    wire [7:0] \AES.r2.t2.t3.in ;
    wire [31:0] \AES.r2.t2.t3.out ;
    wire [7:0] \AES.r2.t2.t3.k0 ;
    wire [7:0] \AES.r2.t2.t3.k1 ;
    wire \AES.r2.t2.t3.s0.clk ;
    wire [7:0] \AES.r2.t2.t3.s0.in ;
    reg [7:0] \AES.r2.t2.t3.s0.out ;
    wire \AES.r2.t2.t3.s4.clk ;
    wire [7:0] \AES.r2.t2.t3.s4.in ;
    reg [7:0] \AES.r2.t2.t3.s4.out ;
    wire \AES.r2.t3.clk ;
    wire [31:0] \AES.r2.t3.state ;
    wire [31:0] \AES.r2.t3.p0 ;
    wire [31:0] \AES.r2.t3.p1 ;
    wire [31:0] \AES.r2.t3.p2 ;
    wire [31:0] \AES.r2.t3.p3 ;
    wire [7:0] \AES.r2.t3.b0 ;
    wire [7:0] \AES.r2.t3.b1 ;
    wire [7:0] \AES.r2.t3.b2 ;
    wire [7:0] \AES.r2.t3.b3 ;
    wire [31:0] \AES.r2.t3.k0 ;
    wire [31:0] \AES.r2.t3.k1 ;
    wire [31:0] \AES.r2.t3.k2 ;
    wire \AES.r2.t3.t0.clk ;
    wire [7:0] \AES.r2.t3.t0.in ;
    wire [31:0] \AES.r2.t3.t0.out ;
    wire [7:0] \AES.r2.t3.t0.k0 ;
    wire [7:0] \AES.r2.t3.t0.k1 ;
    wire \AES.r2.t3.t0.s0.clk ;
    wire [7:0] \AES.r2.t3.t0.s0.in ;
    reg [7:0] \AES.r2.t3.t0.s0.out ;
    wire \AES.r2.t3.t0.s4.clk ;
    wire [7:0] \AES.r2.t3.t0.s4.in ;
    reg [7:0] \AES.r2.t3.t0.s4.out ;
    wire \AES.r2.t3.t1.clk ;
    wire [7:0] \AES.r2.t3.t1.in ;
    wire [31:0] \AES.r2.t3.t1.out ;
    wire [7:0] \AES.r2.t3.t1.k0 ;
    wire [7:0] \AES.r2.t3.t1.k1 ;
    wire \AES.r2.t3.t1.s0.clk ;
    wire [7:0] \AES.r2.t3.t1.s0.in ;
    reg [7:0] \AES.r2.t3.t1.s0.out ;
    wire \AES.r2.t3.t1.s4.clk ;
    wire [7:0] \AES.r2.t3.t1.s4.in ;
    reg [7:0] \AES.r2.t3.t1.s4.out ;
    wire \AES.r2.t3.t2.clk ;
    wire [7:0] \AES.r2.t3.t2.in ;
    wire [31:0] \AES.r2.t3.t2.out ;
    wire [7:0] \AES.r2.t3.t2.k0 ;
    wire [7:0] \AES.r2.t3.t2.k1 ;
    wire \AES.r2.t3.t2.s0.clk ;
    wire [7:0] \AES.r2.t3.t2.s0.in ;
    reg [7:0] \AES.r2.t3.t2.s0.out ;
    wire \AES.r2.t3.t2.s4.clk ;
    wire [7:0] \AES.r2.t3.t2.s4.in ;
    reg [7:0] \AES.r2.t3.t2.s4.out ;
    wire \AES.r2.t3.t3.clk ;
    wire [7:0] \AES.r2.t3.t3.in ;
    wire [31:0] \AES.r2.t3.t3.out ;
    wire [7:0] \AES.r2.t3.t3.k0 ;
    wire [7:0] \AES.r2.t3.t3.k1 ;
    wire \AES.r2.t3.t3.s0.clk ;
    wire [7:0] \AES.r2.t3.t3.s0.in ;
    reg [7:0] \AES.r2.t3.t3.s0.out ;
    wire \AES.r2.t3.t3.s4.clk ;
    wire [7:0] \AES.r2.t3.t3.s4.in ;
    reg [7:0] \AES.r2.t3.t3.s4.out ;
    wire \AES.r3.clk ;
    wire [127:0] \AES.r3.state_in ;
    wire [127:0] \AES.r3.key ;
    reg [127:0] \AES.r3.state_out ;
    wire [31:0] \AES.r3.s0 ;
    wire [31:0] \AES.r3.s1 ;
    wire [31:0] \AES.r3.s2 ;
    wire [31:0] \AES.r3.s3 ;
    wire [31:0] \AES.r3.z0 ;
    wire [31:0] \AES.r3.z1 ;
    wire [31:0] \AES.r3.z2 ;
    wire [31:0] \AES.r3.z3 ;
    wire [31:0] \AES.r3.p00 ;
    wire [31:0] \AES.r3.p01 ;
    wire [31:0] \AES.r3.p02 ;
    wire [31:0] \AES.r3.p03 ;
    wire [31:0] \AES.r3.p10 ;
    wire [31:0] \AES.r3.p11 ;
    wire [31:0] \AES.r3.p12 ;
    wire [31:0] \AES.r3.p13 ;
    wire [31:0] \AES.r3.p20 ;
    wire [31:0] \AES.r3.p21 ;
    wire [31:0] \AES.r3.p22 ;
    wire [31:0] \AES.r3.p23 ;
    wire [31:0] \AES.r3.p30 ;
    wire [31:0] \AES.r3.p31 ;
    wire [31:0] \AES.r3.p32 ;
    wire [31:0] \AES.r3.p33 ;
    wire [31:0] \AES.r3.k0 ;
    wire [31:0] \AES.r3.k1 ;
    wire [31:0] \AES.r3.k2 ;
    wire [31:0] \AES.r3.k3 ;
    wire \AES.r3.t0.clk ;
    wire [31:0] \AES.r3.t0.state ;
    wire [31:0] \AES.r3.t0.p0 ;
    wire [31:0] \AES.r3.t0.p1 ;
    wire [31:0] \AES.r3.t0.p2 ;
    wire [31:0] \AES.r3.t0.p3 ;
    wire [7:0] \AES.r3.t0.b0 ;
    wire [7:0] \AES.r3.t0.b1 ;
    wire [7:0] \AES.r3.t0.b2 ;
    wire [7:0] \AES.r3.t0.b3 ;
    wire [31:0] \AES.r3.t0.k0 ;
    wire [31:0] \AES.r3.t0.k1 ;
    wire [31:0] \AES.r3.t0.k2 ;
    wire \AES.r3.t0.t0.clk ;
    wire [7:0] \AES.r3.t0.t0.in ;
    wire [31:0] \AES.r3.t0.t0.out ;
    wire [7:0] \AES.r3.t0.t0.k0 ;
    wire [7:0] \AES.r3.t0.t0.k1 ;
    wire \AES.r3.t0.t0.s0.clk ;
    wire [7:0] \AES.r3.t0.t0.s0.in ;
    reg [7:0] \AES.r3.t0.t0.s0.out ;
    wire \AES.r3.t0.t0.s4.clk ;
    wire [7:0] \AES.r3.t0.t0.s4.in ;
    reg [7:0] \AES.r3.t0.t0.s4.out ;
    wire \AES.r3.t0.t1.clk ;
    wire [7:0] \AES.r3.t0.t1.in ;
    wire [31:0] \AES.r3.t0.t1.out ;
    wire [7:0] \AES.r3.t0.t1.k0 ;
    wire [7:0] \AES.r3.t0.t1.k1 ;
    wire \AES.r3.t0.t1.s0.clk ;
    wire [7:0] \AES.r3.t0.t1.s0.in ;
    reg [7:0] \AES.r3.t0.t1.s0.out ;
    wire \AES.r3.t0.t1.s4.clk ;
    wire [7:0] \AES.r3.t0.t1.s4.in ;
    reg [7:0] \AES.r3.t0.t1.s4.out ;
    wire \AES.r3.t0.t2.clk ;
    wire [7:0] \AES.r3.t0.t2.in ;
    wire [31:0] \AES.r3.t0.t2.out ;
    wire [7:0] \AES.r3.t0.t2.k0 ;
    wire [7:0] \AES.r3.t0.t2.k1 ;
    wire \AES.r3.t0.t2.s0.clk ;
    wire [7:0] \AES.r3.t0.t2.s0.in ;
    reg [7:0] \AES.r3.t0.t2.s0.out ;
    wire \AES.r3.t0.t2.s4.clk ;
    wire [7:0] \AES.r3.t0.t2.s4.in ;
    reg [7:0] \AES.r3.t0.t2.s4.out ;
    wire \AES.r3.t0.t3.clk ;
    wire [7:0] \AES.r3.t0.t3.in ;
    wire [31:0] \AES.r3.t0.t3.out ;
    wire [7:0] \AES.r3.t0.t3.k0 ;
    wire [7:0] \AES.r3.t0.t3.k1 ;
    wire \AES.r3.t0.t3.s0.clk ;
    wire [7:0] \AES.r3.t0.t3.s0.in ;
    reg [7:0] \AES.r3.t0.t3.s0.out ;
    wire \AES.r3.t0.t3.s4.clk ;
    wire [7:0] \AES.r3.t0.t3.s4.in ;
    reg [7:0] \AES.r3.t0.t3.s4.out ;
    wire \AES.r3.t1.clk ;
    wire [31:0] \AES.r3.t1.state ;
    wire [31:0] \AES.r3.t1.p0 ;
    wire [31:0] \AES.r3.t1.p1 ;
    wire [31:0] \AES.r3.t1.p2 ;
    wire [31:0] \AES.r3.t1.p3 ;
    wire [7:0] \AES.r3.t1.b0 ;
    wire [7:0] \AES.r3.t1.b1 ;
    wire [7:0] \AES.r3.t1.b2 ;
    wire [7:0] \AES.r3.t1.b3 ;
    wire [31:0] \AES.r3.t1.k0 ;
    wire [31:0] \AES.r3.t1.k1 ;
    wire [31:0] \AES.r3.t1.k2 ;
    wire \AES.r3.t1.t0.clk ;
    wire [7:0] \AES.r3.t1.t0.in ;
    wire [31:0] \AES.r3.t1.t0.out ;
    wire [7:0] \AES.r3.t1.t0.k0 ;
    wire [7:0] \AES.r3.t1.t0.k1 ;
    wire \AES.r3.t1.t0.s0.clk ;
    wire [7:0] \AES.r3.t1.t0.s0.in ;
    reg [7:0] \AES.r3.t1.t0.s0.out ;
    wire \AES.r3.t1.t0.s4.clk ;
    wire [7:0] \AES.r3.t1.t0.s4.in ;
    reg [7:0] \AES.r3.t1.t0.s4.out ;
    wire \AES.r3.t1.t1.clk ;
    wire [7:0] \AES.r3.t1.t1.in ;
    wire [31:0] \AES.r3.t1.t1.out ;
    wire [7:0] \AES.r3.t1.t1.k0 ;
    wire [7:0] \AES.r3.t1.t1.k1 ;
    wire \AES.r3.t1.t1.s0.clk ;
    wire [7:0] \AES.r3.t1.t1.s0.in ;
    reg [7:0] \AES.r3.t1.t1.s0.out ;
    wire \AES.r3.t1.t1.s4.clk ;
    wire [7:0] \AES.r3.t1.t1.s4.in ;
    reg [7:0] \AES.r3.t1.t1.s4.out ;
    wire \AES.r3.t1.t2.clk ;
    wire [7:0] \AES.r3.t1.t2.in ;
    wire [31:0] \AES.r3.t1.t2.out ;
    wire [7:0] \AES.r3.t1.t2.k0 ;
    wire [7:0] \AES.r3.t1.t2.k1 ;
    wire \AES.r3.t1.t2.s0.clk ;
    wire [7:0] \AES.r3.t1.t2.s0.in ;
    reg [7:0] \AES.r3.t1.t2.s0.out ;
    wire \AES.r3.t1.t2.s4.clk ;
    wire [7:0] \AES.r3.t1.t2.s4.in ;
    reg [7:0] \AES.r3.t1.t2.s4.out ;
    wire \AES.r3.t1.t3.clk ;
    wire [7:0] \AES.r3.t1.t3.in ;
    wire [31:0] \AES.r3.t1.t3.out ;
    wire [7:0] \AES.r3.t1.t3.k0 ;
    wire [7:0] \AES.r3.t1.t3.k1 ;
    wire \AES.r3.t1.t3.s0.clk ;
    wire [7:0] \AES.r3.t1.t3.s0.in ;
    reg [7:0] \AES.r3.t1.t3.s0.out ;
    wire \AES.r3.t1.t3.s4.clk ;
    wire [7:0] \AES.r3.t1.t3.s4.in ;
    reg [7:0] \AES.r3.t1.t3.s4.out ;
    wire \AES.r3.t2.clk ;
    wire [31:0] \AES.r3.t2.state ;
    wire [31:0] \AES.r3.t2.p0 ;
    wire [31:0] \AES.r3.t2.p1 ;
    wire [31:0] \AES.r3.t2.p2 ;
    wire [31:0] \AES.r3.t2.p3 ;
    wire [7:0] \AES.r3.t2.b0 ;
    wire [7:0] \AES.r3.t2.b1 ;
    wire [7:0] \AES.r3.t2.b2 ;
    wire [7:0] \AES.r3.t2.b3 ;
    wire [31:0] \AES.r3.t2.k0 ;
    wire [31:0] \AES.r3.t2.k1 ;
    wire [31:0] \AES.r3.t2.k2 ;
    wire \AES.r3.t2.t0.clk ;
    wire [7:0] \AES.r3.t2.t0.in ;
    wire [31:0] \AES.r3.t2.t0.out ;
    wire [7:0] \AES.r3.t2.t0.k0 ;
    wire [7:0] \AES.r3.t2.t0.k1 ;
    wire \AES.r3.t2.t0.s0.clk ;
    wire [7:0] \AES.r3.t2.t0.s0.in ;
    reg [7:0] \AES.r3.t2.t0.s0.out ;
    wire \AES.r3.t2.t0.s4.clk ;
    wire [7:0] \AES.r3.t2.t0.s4.in ;
    reg [7:0] \AES.r3.t2.t0.s4.out ;
    wire \AES.r3.t2.t1.clk ;
    wire [7:0] \AES.r3.t2.t1.in ;
    wire [31:0] \AES.r3.t2.t1.out ;
    wire [7:0] \AES.r3.t2.t1.k0 ;
    wire [7:0] \AES.r3.t2.t1.k1 ;
    wire \AES.r3.t2.t1.s0.clk ;
    wire [7:0] \AES.r3.t2.t1.s0.in ;
    reg [7:0] \AES.r3.t2.t1.s0.out ;
    wire \AES.r3.t2.t1.s4.clk ;
    wire [7:0] \AES.r3.t2.t1.s4.in ;
    reg [7:0] \AES.r3.t2.t1.s4.out ;
    wire \AES.r3.t2.t2.clk ;
    wire [7:0] \AES.r3.t2.t2.in ;
    wire [31:0] \AES.r3.t2.t2.out ;
    wire [7:0] \AES.r3.t2.t2.k0 ;
    wire [7:0] \AES.r3.t2.t2.k1 ;
    wire \AES.r3.t2.t2.s0.clk ;
    wire [7:0] \AES.r3.t2.t2.s0.in ;
    reg [7:0] \AES.r3.t2.t2.s0.out ;
    wire \AES.r3.t2.t2.s4.clk ;
    wire [7:0] \AES.r3.t2.t2.s4.in ;
    reg [7:0] \AES.r3.t2.t2.s4.out ;
    wire \AES.r3.t2.t3.clk ;
    wire [7:0] \AES.r3.t2.t3.in ;
    wire [31:0] \AES.r3.t2.t3.out ;
    wire [7:0] \AES.r3.t2.t3.k0 ;
    wire [7:0] \AES.r3.t2.t3.k1 ;
    wire \AES.r3.t2.t3.s0.clk ;
    wire [7:0] \AES.r3.t2.t3.s0.in ;
    reg [7:0] \AES.r3.t2.t3.s0.out ;
    wire \AES.r3.t2.t3.s4.clk ;
    wire [7:0] \AES.r3.t2.t3.s4.in ;
    reg [7:0] \AES.r3.t2.t3.s4.out ;
    wire \AES.r3.t3.clk ;
    wire [31:0] \AES.r3.t3.state ;
    wire [31:0] \AES.r3.t3.p0 ;
    wire [31:0] \AES.r3.t3.p1 ;
    wire [31:0] \AES.r3.t3.p2 ;
    wire [31:0] \AES.r3.t3.p3 ;
    wire [7:0] \AES.r3.t3.b0 ;
    wire [7:0] \AES.r3.t3.b1 ;
    wire [7:0] \AES.r3.t3.b2 ;
    wire [7:0] \AES.r3.t3.b3 ;
    wire [31:0] \AES.r3.t3.k0 ;
    wire [31:0] \AES.r3.t3.k1 ;
    wire [31:0] \AES.r3.t3.k2 ;
    wire \AES.r3.t3.t0.clk ;
    wire [7:0] \AES.r3.t3.t0.in ;
    wire [31:0] \AES.r3.t3.t0.out ;
    wire [7:0] \AES.r3.t3.t0.k0 ;
    wire [7:0] \AES.r3.t3.t0.k1 ;
    wire \AES.r3.t3.t0.s0.clk ;
    wire [7:0] \AES.r3.t3.t0.s0.in ;
    reg [7:0] \AES.r3.t3.t0.s0.out ;
    wire \AES.r3.t3.t0.s4.clk ;
    wire [7:0] \AES.r3.t3.t0.s4.in ;
    reg [7:0] \AES.r3.t3.t0.s4.out ;
    wire \AES.r3.t3.t1.clk ;
    wire [7:0] \AES.r3.t3.t1.in ;
    wire [31:0] \AES.r3.t3.t1.out ;
    wire [7:0] \AES.r3.t3.t1.k0 ;
    wire [7:0] \AES.r3.t3.t1.k1 ;
    wire \AES.r3.t3.t1.s0.clk ;
    wire [7:0] \AES.r3.t3.t1.s0.in ;
    reg [7:0] \AES.r3.t3.t1.s0.out ;
    wire \AES.r3.t3.t1.s4.clk ;
    wire [7:0] \AES.r3.t3.t1.s4.in ;
    reg [7:0] \AES.r3.t3.t1.s4.out ;
    wire \AES.r3.t3.t2.clk ;
    wire [7:0] \AES.r3.t3.t2.in ;
    wire [31:0] \AES.r3.t3.t2.out ;
    wire [7:0] \AES.r3.t3.t2.k0 ;
    wire [7:0] \AES.r3.t3.t2.k1 ;
    wire \AES.r3.t3.t2.s0.clk ;
    wire [7:0] \AES.r3.t3.t2.s0.in ;
    reg [7:0] \AES.r3.t3.t2.s0.out ;
    wire \AES.r3.t3.t2.s4.clk ;
    wire [7:0] \AES.r3.t3.t2.s4.in ;
    reg [7:0] \AES.r3.t3.t2.s4.out ;
    wire \AES.r3.t3.t3.clk ;
    wire [7:0] \AES.r3.t3.t3.in ;
    wire [31:0] \AES.r3.t3.t3.out ;
    wire [7:0] \AES.r3.t3.t3.k0 ;
    wire [7:0] \AES.r3.t3.t3.k1 ;
    wire \AES.r3.t3.t3.s0.clk ;
    wire [7:0] \AES.r3.t3.t3.s0.in ;
    reg [7:0] \AES.r3.t3.t3.s0.out ;
    wire \AES.r3.t3.t3.s4.clk ;
    wire [7:0] \AES.r3.t3.t3.s4.in ;
    reg [7:0] \AES.r3.t3.t3.s4.out ;
    wire \AES.r4.clk ;
    wire [127:0] \AES.r4.state_in ;
    wire [127:0] \AES.r4.key ;
    reg [127:0] \AES.r4.state_out ;
    wire [31:0] \AES.r4.s0 ;
    wire [31:0] \AES.r4.s1 ;
    wire [31:0] \AES.r4.s2 ;
    wire [31:0] \AES.r4.s3 ;
    wire [31:0] \AES.r4.z0 ;
    wire [31:0] \AES.r4.z1 ;
    wire [31:0] \AES.r4.z2 ;
    wire [31:0] \AES.r4.z3 ;
    wire [31:0] \AES.r4.p00 ;
    wire [31:0] \AES.r4.p01 ;
    wire [31:0] \AES.r4.p02 ;
    wire [31:0] \AES.r4.p03 ;
    wire [31:0] \AES.r4.p10 ;
    wire [31:0] \AES.r4.p11 ;
    wire [31:0] \AES.r4.p12 ;
    wire [31:0] \AES.r4.p13 ;
    wire [31:0] \AES.r4.p20 ;
    wire [31:0] \AES.r4.p21 ;
    wire [31:0] \AES.r4.p22 ;
    wire [31:0] \AES.r4.p23 ;
    wire [31:0] \AES.r4.p30 ;
    wire [31:0] \AES.r4.p31 ;
    wire [31:0] \AES.r4.p32 ;
    wire [31:0] \AES.r4.p33 ;
    wire [31:0] \AES.r4.k0 ;
    wire [31:0] \AES.r4.k1 ;
    wire [31:0] \AES.r4.k2 ;
    wire [31:0] \AES.r4.k3 ;
    wire \AES.r4.t0.clk ;
    wire [31:0] \AES.r4.t0.state ;
    wire [31:0] \AES.r4.t0.p0 ;
    wire [31:0] \AES.r4.t0.p1 ;
    wire [31:0] \AES.r4.t0.p2 ;
    wire [31:0] \AES.r4.t0.p3 ;
    wire [7:0] \AES.r4.t0.b0 ;
    wire [7:0] \AES.r4.t0.b1 ;
    wire [7:0] \AES.r4.t0.b2 ;
    wire [7:0] \AES.r4.t0.b3 ;
    wire [31:0] \AES.r4.t0.k0 ;
    wire [31:0] \AES.r4.t0.k1 ;
    wire [31:0] \AES.r4.t0.k2 ;
    wire \AES.r4.t0.t0.clk ;
    wire [7:0] \AES.r4.t0.t0.in ;
    wire [31:0] \AES.r4.t0.t0.out ;
    wire [7:0] \AES.r4.t0.t0.k0 ;
    wire [7:0] \AES.r4.t0.t0.k1 ;
    wire \AES.r4.t0.t0.s0.clk ;
    wire [7:0] \AES.r4.t0.t0.s0.in ;
    reg [7:0] \AES.r4.t0.t0.s0.out ;
    wire \AES.r4.t0.t0.s4.clk ;
    wire [7:0] \AES.r4.t0.t0.s4.in ;
    reg [7:0] \AES.r4.t0.t0.s4.out ;
    wire \AES.r4.t0.t1.clk ;
    wire [7:0] \AES.r4.t0.t1.in ;
    wire [31:0] \AES.r4.t0.t1.out ;
    wire [7:0] \AES.r4.t0.t1.k0 ;
    wire [7:0] \AES.r4.t0.t1.k1 ;
    wire \AES.r4.t0.t1.s0.clk ;
    wire [7:0] \AES.r4.t0.t1.s0.in ;
    reg [7:0] \AES.r4.t0.t1.s0.out ;
    wire \AES.r4.t0.t1.s4.clk ;
    wire [7:0] \AES.r4.t0.t1.s4.in ;
    reg [7:0] \AES.r4.t0.t1.s4.out ;
    wire \AES.r4.t0.t2.clk ;
    wire [7:0] \AES.r4.t0.t2.in ;
    wire [31:0] \AES.r4.t0.t2.out ;
    wire [7:0] \AES.r4.t0.t2.k0 ;
    wire [7:0] \AES.r4.t0.t2.k1 ;
    wire \AES.r4.t0.t2.s0.clk ;
    wire [7:0] \AES.r4.t0.t2.s0.in ;
    reg [7:0] \AES.r4.t0.t2.s0.out ;
    wire \AES.r4.t0.t2.s4.clk ;
    wire [7:0] \AES.r4.t0.t2.s4.in ;
    reg [7:0] \AES.r4.t0.t2.s4.out ;
    wire \AES.r4.t0.t3.clk ;
    wire [7:0] \AES.r4.t0.t3.in ;
    wire [31:0] \AES.r4.t0.t3.out ;
    wire [7:0] \AES.r4.t0.t3.k0 ;
    wire [7:0] \AES.r4.t0.t3.k1 ;
    wire \AES.r4.t0.t3.s0.clk ;
    wire [7:0] \AES.r4.t0.t3.s0.in ;
    reg [7:0] \AES.r4.t0.t3.s0.out ;
    wire \AES.r4.t0.t3.s4.clk ;
    wire [7:0] \AES.r4.t0.t3.s4.in ;
    reg [7:0] \AES.r4.t0.t3.s4.out ;
    wire \AES.r4.t1.clk ;
    wire [31:0] \AES.r4.t1.state ;
    wire [31:0] \AES.r4.t1.p0 ;
    wire [31:0] \AES.r4.t1.p1 ;
    wire [31:0] \AES.r4.t1.p2 ;
    wire [31:0] \AES.r4.t1.p3 ;
    wire [7:0] \AES.r4.t1.b0 ;
    wire [7:0] \AES.r4.t1.b1 ;
    wire [7:0] \AES.r4.t1.b2 ;
    wire [7:0] \AES.r4.t1.b3 ;
    wire [31:0] \AES.r4.t1.k0 ;
    wire [31:0] \AES.r4.t1.k1 ;
    wire [31:0] \AES.r4.t1.k2 ;
    wire \AES.r4.t1.t0.clk ;
    wire [7:0] \AES.r4.t1.t0.in ;
    wire [31:0] \AES.r4.t1.t0.out ;
    wire [7:0] \AES.r4.t1.t0.k0 ;
    wire [7:0] \AES.r4.t1.t0.k1 ;
    wire \AES.r4.t1.t0.s0.clk ;
    wire [7:0] \AES.r4.t1.t0.s0.in ;
    reg [7:0] \AES.r4.t1.t0.s0.out ;
    wire \AES.r4.t1.t0.s4.clk ;
    wire [7:0] \AES.r4.t1.t0.s4.in ;
    reg [7:0] \AES.r4.t1.t0.s4.out ;
    wire \AES.r4.t1.t1.clk ;
    wire [7:0] \AES.r4.t1.t1.in ;
    wire [31:0] \AES.r4.t1.t1.out ;
    wire [7:0] \AES.r4.t1.t1.k0 ;
    wire [7:0] \AES.r4.t1.t1.k1 ;
    wire \AES.r4.t1.t1.s0.clk ;
    wire [7:0] \AES.r4.t1.t1.s0.in ;
    reg [7:0] \AES.r4.t1.t1.s0.out ;
    wire \AES.r4.t1.t1.s4.clk ;
    wire [7:0] \AES.r4.t1.t1.s4.in ;
    reg [7:0] \AES.r4.t1.t1.s4.out ;
    wire \AES.r4.t1.t2.clk ;
    wire [7:0] \AES.r4.t1.t2.in ;
    wire [31:0] \AES.r4.t1.t2.out ;
    wire [7:0] \AES.r4.t1.t2.k0 ;
    wire [7:0] \AES.r4.t1.t2.k1 ;
    wire \AES.r4.t1.t2.s0.clk ;
    wire [7:0] \AES.r4.t1.t2.s0.in ;
    reg [7:0] \AES.r4.t1.t2.s0.out ;
    wire \AES.r4.t1.t2.s4.clk ;
    wire [7:0] \AES.r4.t1.t2.s4.in ;
    reg [7:0] \AES.r4.t1.t2.s4.out ;
    wire \AES.r4.t1.t3.clk ;
    wire [7:0] \AES.r4.t1.t3.in ;
    wire [31:0] \AES.r4.t1.t3.out ;
    wire [7:0] \AES.r4.t1.t3.k0 ;
    wire [7:0] \AES.r4.t1.t3.k1 ;
    wire \AES.r4.t1.t3.s0.clk ;
    wire [7:0] \AES.r4.t1.t3.s0.in ;
    reg [7:0] \AES.r4.t1.t3.s0.out ;
    wire \AES.r4.t1.t3.s4.clk ;
    wire [7:0] \AES.r4.t1.t3.s4.in ;
    reg [7:0] \AES.r4.t1.t3.s4.out ;
    wire \AES.r4.t2.clk ;
    wire [31:0] \AES.r4.t2.state ;
    wire [31:0] \AES.r4.t2.p0 ;
    wire [31:0] \AES.r4.t2.p1 ;
    wire [31:0] \AES.r4.t2.p2 ;
    wire [31:0] \AES.r4.t2.p3 ;
    wire [7:0] \AES.r4.t2.b0 ;
    wire [7:0] \AES.r4.t2.b1 ;
    wire [7:0] \AES.r4.t2.b2 ;
    wire [7:0] \AES.r4.t2.b3 ;
    wire [31:0] \AES.r4.t2.k0 ;
    wire [31:0] \AES.r4.t2.k1 ;
    wire [31:0] \AES.r4.t2.k2 ;
    wire \AES.r4.t2.t0.clk ;
    wire [7:0] \AES.r4.t2.t0.in ;
    wire [31:0] \AES.r4.t2.t0.out ;
    wire [7:0] \AES.r4.t2.t0.k0 ;
    wire [7:0] \AES.r4.t2.t0.k1 ;
    wire \AES.r4.t2.t0.s0.clk ;
    wire [7:0] \AES.r4.t2.t0.s0.in ;
    reg [7:0] \AES.r4.t2.t0.s0.out ;
    wire \AES.r4.t2.t0.s4.clk ;
    wire [7:0] \AES.r4.t2.t0.s4.in ;
    reg [7:0] \AES.r4.t2.t0.s4.out ;
    wire \AES.r4.t2.t1.clk ;
    wire [7:0] \AES.r4.t2.t1.in ;
    wire [31:0] \AES.r4.t2.t1.out ;
    wire [7:0] \AES.r4.t2.t1.k0 ;
    wire [7:0] \AES.r4.t2.t1.k1 ;
    wire \AES.r4.t2.t1.s0.clk ;
    wire [7:0] \AES.r4.t2.t1.s0.in ;
    reg [7:0] \AES.r4.t2.t1.s0.out ;
    wire \AES.r4.t2.t1.s4.clk ;
    wire [7:0] \AES.r4.t2.t1.s4.in ;
    reg [7:0] \AES.r4.t2.t1.s4.out ;
    wire \AES.r4.t2.t2.clk ;
    wire [7:0] \AES.r4.t2.t2.in ;
    wire [31:0] \AES.r4.t2.t2.out ;
    wire [7:0] \AES.r4.t2.t2.k0 ;
    wire [7:0] \AES.r4.t2.t2.k1 ;
    wire \AES.r4.t2.t2.s0.clk ;
    wire [7:0] \AES.r4.t2.t2.s0.in ;
    reg [7:0] \AES.r4.t2.t2.s0.out ;
    wire \AES.r4.t2.t2.s4.clk ;
    wire [7:0] \AES.r4.t2.t2.s4.in ;
    reg [7:0] \AES.r4.t2.t2.s4.out ;
    wire \AES.r4.t2.t3.clk ;
    wire [7:0] \AES.r4.t2.t3.in ;
    wire [31:0] \AES.r4.t2.t3.out ;
    wire [7:0] \AES.r4.t2.t3.k0 ;
    wire [7:0] \AES.r4.t2.t3.k1 ;
    wire \AES.r4.t2.t3.s0.clk ;
    wire [7:0] \AES.r4.t2.t3.s0.in ;
    reg [7:0] \AES.r4.t2.t3.s0.out ;
    wire \AES.r4.t2.t3.s4.clk ;
    wire [7:0] \AES.r4.t2.t3.s4.in ;
    reg [7:0] \AES.r4.t2.t3.s4.out ;
    wire \AES.r4.t3.clk ;
    wire [31:0] \AES.r4.t3.state ;
    wire [31:0] \AES.r4.t3.p0 ;
    wire [31:0] \AES.r4.t3.p1 ;
    wire [31:0] \AES.r4.t3.p2 ;
    wire [31:0] \AES.r4.t3.p3 ;
    wire [7:0] \AES.r4.t3.b0 ;
    wire [7:0] \AES.r4.t3.b1 ;
    wire [7:0] \AES.r4.t3.b2 ;
    wire [7:0] \AES.r4.t3.b3 ;
    wire [31:0] \AES.r4.t3.k0 ;
    wire [31:0] \AES.r4.t3.k1 ;
    wire [31:0] \AES.r4.t3.k2 ;
    wire \AES.r4.t3.t0.clk ;
    wire [7:0] \AES.r4.t3.t0.in ;
    wire [31:0] \AES.r4.t3.t0.out ;
    wire [7:0] \AES.r4.t3.t0.k0 ;
    wire [7:0] \AES.r4.t3.t0.k1 ;
    wire \AES.r4.t3.t0.s0.clk ;
    wire [7:0] \AES.r4.t3.t0.s0.in ;
    reg [7:0] \AES.r4.t3.t0.s0.out ;
    wire \AES.r4.t3.t0.s4.clk ;
    wire [7:0] \AES.r4.t3.t0.s4.in ;
    reg [7:0] \AES.r4.t3.t0.s4.out ;
    wire \AES.r4.t3.t1.clk ;
    wire [7:0] \AES.r4.t3.t1.in ;
    wire [31:0] \AES.r4.t3.t1.out ;
    wire [7:0] \AES.r4.t3.t1.k0 ;
    wire [7:0] \AES.r4.t3.t1.k1 ;
    wire \AES.r4.t3.t1.s0.clk ;
    wire [7:0] \AES.r4.t3.t1.s0.in ;
    reg [7:0] \AES.r4.t3.t1.s0.out ;
    wire \AES.r4.t3.t1.s4.clk ;
    wire [7:0] \AES.r4.t3.t1.s4.in ;
    reg [7:0] \AES.r4.t3.t1.s4.out ;
    wire \AES.r4.t3.t2.clk ;
    wire [7:0] \AES.r4.t3.t2.in ;
    wire [31:0] \AES.r4.t3.t2.out ;
    wire [7:0] \AES.r4.t3.t2.k0 ;
    wire [7:0] \AES.r4.t3.t2.k1 ;
    wire \AES.r4.t3.t2.s0.clk ;
    wire [7:0] \AES.r4.t3.t2.s0.in ;
    reg [7:0] \AES.r4.t3.t2.s0.out ;
    wire \AES.r4.t3.t2.s4.clk ;
    wire [7:0] \AES.r4.t3.t2.s4.in ;
    reg [7:0] \AES.r4.t3.t2.s4.out ;
    wire \AES.r4.t3.t3.clk ;
    wire [7:0] \AES.r4.t3.t3.in ;
    wire [31:0] \AES.r4.t3.t3.out ;
    wire [7:0] \AES.r4.t3.t3.k0 ;
    wire [7:0] \AES.r4.t3.t3.k1 ;
    wire \AES.r4.t3.t3.s0.clk ;
    wire [7:0] \AES.r4.t3.t3.s0.in ;
    reg [7:0] \AES.r4.t3.t3.s0.out ;
    wire \AES.r4.t3.t3.s4.clk ;
    wire [7:0] \AES.r4.t3.t3.s4.in ;
    reg [7:0] \AES.r4.t3.t3.s4.out ;
    wire \AES.r5.clk ;
    wire [127:0] \AES.r5.state_in ;
    wire [127:0] \AES.r5.key ;
    reg [127:0] \AES.r5.state_out ;
    wire [31:0] \AES.r5.s0 ;
    wire [31:0] \AES.r5.s1 ;
    wire [31:0] \AES.r5.s2 ;
    wire [31:0] \AES.r5.s3 ;
    wire [31:0] \AES.r5.z0 ;
    wire [31:0] \AES.r5.z1 ;
    wire [31:0] \AES.r5.z2 ;
    wire [31:0] \AES.r5.z3 ;
    wire [31:0] \AES.r5.p00 ;
    wire [31:0] \AES.r5.p01 ;
    wire [31:0] \AES.r5.p02 ;
    wire [31:0] \AES.r5.p03 ;
    wire [31:0] \AES.r5.p10 ;
    wire [31:0] \AES.r5.p11 ;
    wire [31:0] \AES.r5.p12 ;
    wire [31:0] \AES.r5.p13 ;
    wire [31:0] \AES.r5.p20 ;
    wire [31:0] \AES.r5.p21 ;
    wire [31:0] \AES.r5.p22 ;
    wire [31:0] \AES.r5.p23 ;
    wire [31:0] \AES.r5.p30 ;
    wire [31:0] \AES.r5.p31 ;
    wire [31:0] \AES.r5.p32 ;
    wire [31:0] \AES.r5.p33 ;
    wire [31:0] \AES.r5.k0 ;
    wire [31:0] \AES.r5.k1 ;
    wire [31:0] \AES.r5.k2 ;
    wire [31:0] \AES.r5.k3 ;
    wire \AES.r5.t0.clk ;
    wire [31:0] \AES.r5.t0.state ;
    wire [31:0] \AES.r5.t0.p0 ;
    wire [31:0] \AES.r5.t0.p1 ;
    wire [31:0] \AES.r5.t0.p2 ;
    wire [31:0] \AES.r5.t0.p3 ;
    wire [7:0] \AES.r5.t0.b0 ;
    wire [7:0] \AES.r5.t0.b1 ;
    wire [7:0] \AES.r5.t0.b2 ;
    wire [7:0] \AES.r5.t0.b3 ;
    wire [31:0] \AES.r5.t0.k0 ;
    wire [31:0] \AES.r5.t0.k1 ;
    wire [31:0] \AES.r5.t0.k2 ;
    wire \AES.r5.t0.t0.clk ;
    wire [7:0] \AES.r5.t0.t0.in ;
    wire [31:0] \AES.r5.t0.t0.out ;
    wire [7:0] \AES.r5.t0.t0.k0 ;
    wire [7:0] \AES.r5.t0.t0.k1 ;
    wire \AES.r5.t0.t0.s0.clk ;
    wire [7:0] \AES.r5.t0.t0.s0.in ;
    reg [7:0] \AES.r5.t0.t0.s0.out ;
    wire \AES.r5.t0.t0.s4.clk ;
    wire [7:0] \AES.r5.t0.t0.s4.in ;
    reg [7:0] \AES.r5.t0.t0.s4.out ;
    wire \AES.r5.t0.t1.clk ;
    wire [7:0] \AES.r5.t0.t1.in ;
    wire [31:0] \AES.r5.t0.t1.out ;
    wire [7:0] \AES.r5.t0.t1.k0 ;
    wire [7:0] \AES.r5.t0.t1.k1 ;
    wire \AES.r5.t0.t1.s0.clk ;
    wire [7:0] \AES.r5.t0.t1.s0.in ;
    reg [7:0] \AES.r5.t0.t1.s0.out ;
    wire \AES.r5.t0.t1.s4.clk ;
    wire [7:0] \AES.r5.t0.t1.s4.in ;
    reg [7:0] \AES.r5.t0.t1.s4.out ;
    wire \AES.r5.t0.t2.clk ;
    wire [7:0] \AES.r5.t0.t2.in ;
    wire [31:0] \AES.r5.t0.t2.out ;
    wire [7:0] \AES.r5.t0.t2.k0 ;
    wire [7:0] \AES.r5.t0.t2.k1 ;
    wire \AES.r5.t0.t2.s0.clk ;
    wire [7:0] \AES.r5.t0.t2.s0.in ;
    reg [7:0] \AES.r5.t0.t2.s0.out ;
    wire \AES.r5.t0.t2.s4.clk ;
    wire [7:0] \AES.r5.t0.t2.s4.in ;
    reg [7:0] \AES.r5.t0.t2.s4.out ;
    wire \AES.r5.t0.t3.clk ;
    wire [7:0] \AES.r5.t0.t3.in ;
    wire [31:0] \AES.r5.t0.t3.out ;
    wire [7:0] \AES.r5.t0.t3.k0 ;
    wire [7:0] \AES.r5.t0.t3.k1 ;
    wire \AES.r5.t0.t3.s0.clk ;
    wire [7:0] \AES.r5.t0.t3.s0.in ;
    reg [7:0] \AES.r5.t0.t3.s0.out ;
    wire \AES.r5.t0.t3.s4.clk ;
    wire [7:0] \AES.r5.t0.t3.s4.in ;
    reg [7:0] \AES.r5.t0.t3.s4.out ;
    wire \AES.r5.t1.clk ;
    wire [31:0] \AES.r5.t1.state ;
    wire [31:0] \AES.r5.t1.p0 ;
    wire [31:0] \AES.r5.t1.p1 ;
    wire [31:0] \AES.r5.t1.p2 ;
    wire [31:0] \AES.r5.t1.p3 ;
    wire [7:0] \AES.r5.t1.b0 ;
    wire [7:0] \AES.r5.t1.b1 ;
    wire [7:0] \AES.r5.t1.b2 ;
    wire [7:0] \AES.r5.t1.b3 ;
    wire [31:0] \AES.r5.t1.k0 ;
    wire [31:0] \AES.r5.t1.k1 ;
    wire [31:0] \AES.r5.t1.k2 ;
    wire \AES.r5.t1.t0.clk ;
    wire [7:0] \AES.r5.t1.t0.in ;
    wire [31:0] \AES.r5.t1.t0.out ;
    wire [7:0] \AES.r5.t1.t0.k0 ;
    wire [7:0] \AES.r5.t1.t0.k1 ;
    wire \AES.r5.t1.t0.s0.clk ;
    wire [7:0] \AES.r5.t1.t0.s0.in ;
    reg [7:0] \AES.r5.t1.t0.s0.out ;
    wire \AES.r5.t1.t0.s4.clk ;
    wire [7:0] \AES.r5.t1.t0.s4.in ;
    reg [7:0] \AES.r5.t1.t0.s4.out ;
    wire \AES.r5.t1.t1.clk ;
    wire [7:0] \AES.r5.t1.t1.in ;
    wire [31:0] \AES.r5.t1.t1.out ;
    wire [7:0] \AES.r5.t1.t1.k0 ;
    wire [7:0] \AES.r5.t1.t1.k1 ;
    wire \AES.r5.t1.t1.s0.clk ;
    wire [7:0] \AES.r5.t1.t1.s0.in ;
    reg [7:0] \AES.r5.t1.t1.s0.out ;
    wire \AES.r5.t1.t1.s4.clk ;
    wire [7:0] \AES.r5.t1.t1.s4.in ;
    reg [7:0] \AES.r5.t1.t1.s4.out ;
    wire \AES.r5.t1.t2.clk ;
    wire [7:0] \AES.r5.t1.t2.in ;
    wire [31:0] \AES.r5.t1.t2.out ;
    wire [7:0] \AES.r5.t1.t2.k0 ;
    wire [7:0] \AES.r5.t1.t2.k1 ;
    wire \AES.r5.t1.t2.s0.clk ;
    wire [7:0] \AES.r5.t1.t2.s0.in ;
    reg [7:0] \AES.r5.t1.t2.s0.out ;
    wire \AES.r5.t1.t2.s4.clk ;
    wire [7:0] \AES.r5.t1.t2.s4.in ;
    reg [7:0] \AES.r5.t1.t2.s4.out ;
    wire \AES.r5.t1.t3.clk ;
    wire [7:0] \AES.r5.t1.t3.in ;
    wire [31:0] \AES.r5.t1.t3.out ;
    wire [7:0] \AES.r5.t1.t3.k0 ;
    wire [7:0] \AES.r5.t1.t3.k1 ;
    wire \AES.r5.t1.t3.s0.clk ;
    wire [7:0] \AES.r5.t1.t3.s0.in ;
    reg [7:0] \AES.r5.t1.t3.s0.out ;
    wire \AES.r5.t1.t3.s4.clk ;
    wire [7:0] \AES.r5.t1.t3.s4.in ;
    reg [7:0] \AES.r5.t1.t3.s4.out ;
    wire \AES.r5.t2.clk ;
    wire [31:0] \AES.r5.t2.state ;
    wire [31:0] \AES.r5.t2.p0 ;
    wire [31:0] \AES.r5.t2.p1 ;
    wire [31:0] \AES.r5.t2.p2 ;
    wire [31:0] \AES.r5.t2.p3 ;
    wire [7:0] \AES.r5.t2.b0 ;
    wire [7:0] \AES.r5.t2.b1 ;
    wire [7:0] \AES.r5.t2.b2 ;
    wire [7:0] \AES.r5.t2.b3 ;
    wire [31:0] \AES.r5.t2.k0 ;
    wire [31:0] \AES.r5.t2.k1 ;
    wire [31:0] \AES.r5.t2.k2 ;
    wire \AES.r5.t2.t0.clk ;
    wire [7:0] \AES.r5.t2.t0.in ;
    wire [31:0] \AES.r5.t2.t0.out ;
    wire [7:0] \AES.r5.t2.t0.k0 ;
    wire [7:0] \AES.r5.t2.t0.k1 ;
    wire \AES.r5.t2.t0.s0.clk ;
    wire [7:0] \AES.r5.t2.t0.s0.in ;
    reg [7:0] \AES.r5.t2.t0.s0.out ;
    wire \AES.r5.t2.t0.s4.clk ;
    wire [7:0] \AES.r5.t2.t0.s4.in ;
    reg [7:0] \AES.r5.t2.t0.s4.out ;
    wire \AES.r5.t2.t1.clk ;
    wire [7:0] \AES.r5.t2.t1.in ;
    wire [31:0] \AES.r5.t2.t1.out ;
    wire [7:0] \AES.r5.t2.t1.k0 ;
    wire [7:0] \AES.r5.t2.t1.k1 ;
    wire \AES.r5.t2.t1.s0.clk ;
    wire [7:0] \AES.r5.t2.t1.s0.in ;
    reg [7:0] \AES.r5.t2.t1.s0.out ;
    wire \AES.r5.t2.t1.s4.clk ;
    wire [7:0] \AES.r5.t2.t1.s4.in ;
    reg [7:0] \AES.r5.t2.t1.s4.out ;
    wire \AES.r5.t2.t2.clk ;
    wire [7:0] \AES.r5.t2.t2.in ;
    wire [31:0] \AES.r5.t2.t2.out ;
    wire [7:0] \AES.r5.t2.t2.k0 ;
    wire [7:0] \AES.r5.t2.t2.k1 ;
    wire \AES.r5.t2.t2.s0.clk ;
    wire [7:0] \AES.r5.t2.t2.s0.in ;
    reg [7:0] \AES.r5.t2.t2.s0.out ;
    wire \AES.r5.t2.t2.s4.clk ;
    wire [7:0] \AES.r5.t2.t2.s4.in ;
    reg [7:0] \AES.r5.t2.t2.s4.out ;
    wire \AES.r5.t2.t3.clk ;
    wire [7:0] \AES.r5.t2.t3.in ;
    wire [31:0] \AES.r5.t2.t3.out ;
    wire [7:0] \AES.r5.t2.t3.k0 ;
    wire [7:0] \AES.r5.t2.t3.k1 ;
    wire \AES.r5.t2.t3.s0.clk ;
    wire [7:0] \AES.r5.t2.t3.s0.in ;
    reg [7:0] \AES.r5.t2.t3.s0.out ;
    wire \AES.r5.t2.t3.s4.clk ;
    wire [7:0] \AES.r5.t2.t3.s4.in ;
    reg [7:0] \AES.r5.t2.t3.s4.out ;
    wire \AES.r5.t3.clk ;
    wire [31:0] \AES.r5.t3.state ;
    wire [31:0] \AES.r5.t3.p0 ;
    wire [31:0] \AES.r5.t3.p1 ;
    wire [31:0] \AES.r5.t3.p2 ;
    wire [31:0] \AES.r5.t3.p3 ;
    wire [7:0] \AES.r5.t3.b0 ;
    wire [7:0] \AES.r5.t3.b1 ;
    wire [7:0] \AES.r5.t3.b2 ;
    wire [7:0] \AES.r5.t3.b3 ;
    wire [31:0] \AES.r5.t3.k0 ;
    wire [31:0] \AES.r5.t3.k1 ;
    wire [31:0] \AES.r5.t3.k2 ;
    wire \AES.r5.t3.t0.clk ;
    wire [7:0] \AES.r5.t3.t0.in ;
    wire [31:0] \AES.r5.t3.t0.out ;
    wire [7:0] \AES.r5.t3.t0.k0 ;
    wire [7:0] \AES.r5.t3.t0.k1 ;
    wire \AES.r5.t3.t0.s0.clk ;
    wire [7:0] \AES.r5.t3.t0.s0.in ;
    reg [7:0] \AES.r5.t3.t0.s0.out ;
    wire \AES.r5.t3.t0.s4.clk ;
    wire [7:0] \AES.r5.t3.t0.s4.in ;
    reg [7:0] \AES.r5.t3.t0.s4.out ;
    wire \AES.r5.t3.t1.clk ;
    wire [7:0] \AES.r5.t3.t1.in ;
    wire [31:0] \AES.r5.t3.t1.out ;
    wire [7:0] \AES.r5.t3.t1.k0 ;
    wire [7:0] \AES.r5.t3.t1.k1 ;
    wire \AES.r5.t3.t1.s0.clk ;
    wire [7:0] \AES.r5.t3.t1.s0.in ;
    reg [7:0] \AES.r5.t3.t1.s0.out ;
    wire \AES.r5.t3.t1.s4.clk ;
    wire [7:0] \AES.r5.t3.t1.s4.in ;
    reg [7:0] \AES.r5.t3.t1.s4.out ;
    wire \AES.r5.t3.t2.clk ;
    wire [7:0] \AES.r5.t3.t2.in ;
    wire [31:0] \AES.r5.t3.t2.out ;
    wire [7:0] \AES.r5.t3.t2.k0 ;
    wire [7:0] \AES.r5.t3.t2.k1 ;
    wire \AES.r5.t3.t2.s0.clk ;
    wire [7:0] \AES.r5.t3.t2.s0.in ;
    reg [7:0] \AES.r5.t3.t2.s0.out ;
    wire \AES.r5.t3.t2.s4.clk ;
    wire [7:0] \AES.r5.t3.t2.s4.in ;
    reg [7:0] \AES.r5.t3.t2.s4.out ;
    wire \AES.r5.t3.t3.clk ;
    wire [7:0] \AES.r5.t3.t3.in ;
    wire [31:0] \AES.r5.t3.t3.out ;
    wire [7:0] \AES.r5.t3.t3.k0 ;
    wire [7:0] \AES.r5.t3.t3.k1 ;
    wire \AES.r5.t3.t3.s0.clk ;
    wire [7:0] \AES.r5.t3.t3.s0.in ;
    reg [7:0] \AES.r5.t3.t3.s0.out ;
    wire \AES.r5.t3.t3.s4.clk ;
    wire [7:0] \AES.r5.t3.t3.s4.in ;
    reg [7:0] \AES.r5.t3.t3.s4.out ;
    wire \AES.r6.clk ;
    wire [127:0] \AES.r6.state_in ;
    wire [127:0] \AES.r6.key ;
    reg [127:0] \AES.r6.state_out ;
    wire [31:0] \AES.r6.s0 ;
    wire [31:0] \AES.r6.s1 ;
    wire [31:0] \AES.r6.s2 ;
    wire [31:0] \AES.r6.s3 ;
    wire [31:0] \AES.r6.z0 ;
    wire [31:0] \AES.r6.z1 ;
    wire [31:0] \AES.r6.z2 ;
    wire [31:0] \AES.r6.z3 ;
    wire [31:0] \AES.r6.p00 ;
    wire [31:0] \AES.r6.p01 ;
    wire [31:0] \AES.r6.p02 ;
    wire [31:0] \AES.r6.p03 ;
    wire [31:0] \AES.r6.p10 ;
    wire [31:0] \AES.r6.p11 ;
    wire [31:0] \AES.r6.p12 ;
    wire [31:0] \AES.r6.p13 ;
    wire [31:0] \AES.r6.p20 ;
    wire [31:0] \AES.r6.p21 ;
    wire [31:0] \AES.r6.p22 ;
    wire [31:0] \AES.r6.p23 ;
    wire [31:0] \AES.r6.p30 ;
    wire [31:0] \AES.r6.p31 ;
    wire [31:0] \AES.r6.p32 ;
    wire [31:0] \AES.r6.p33 ;
    wire [31:0] \AES.r6.k0 ;
    wire [31:0] \AES.r6.k1 ;
    wire [31:0] \AES.r6.k2 ;
    wire [31:0] \AES.r6.k3 ;
    wire \AES.r6.t0.clk ;
    wire [31:0] \AES.r6.t0.state ;
    wire [31:0] \AES.r6.t0.p0 ;
    wire [31:0] \AES.r6.t0.p1 ;
    wire [31:0] \AES.r6.t0.p2 ;
    wire [31:0] \AES.r6.t0.p3 ;
    wire [7:0] \AES.r6.t0.b0 ;
    wire [7:0] \AES.r6.t0.b1 ;
    wire [7:0] \AES.r6.t0.b2 ;
    wire [7:0] \AES.r6.t0.b3 ;
    wire [31:0] \AES.r6.t0.k0 ;
    wire [31:0] \AES.r6.t0.k1 ;
    wire [31:0] \AES.r6.t0.k2 ;
    wire \AES.r6.t0.t0.clk ;
    wire [7:0] \AES.r6.t0.t0.in ;
    wire [31:0] \AES.r6.t0.t0.out ;
    wire [7:0] \AES.r6.t0.t0.k0 ;
    wire [7:0] \AES.r6.t0.t0.k1 ;
    wire \AES.r6.t0.t0.s0.clk ;
    wire [7:0] \AES.r6.t0.t0.s0.in ;
    reg [7:0] \AES.r6.t0.t0.s0.out ;
    wire \AES.r6.t0.t0.s4.clk ;
    wire [7:0] \AES.r6.t0.t0.s4.in ;
    reg [7:0] \AES.r6.t0.t0.s4.out ;
    wire \AES.r6.t0.t1.clk ;
    wire [7:0] \AES.r6.t0.t1.in ;
    wire [31:0] \AES.r6.t0.t1.out ;
    wire [7:0] \AES.r6.t0.t1.k0 ;
    wire [7:0] \AES.r6.t0.t1.k1 ;
    wire \AES.r6.t0.t1.s0.clk ;
    wire [7:0] \AES.r6.t0.t1.s0.in ;
    reg [7:0] \AES.r6.t0.t1.s0.out ;
    wire \AES.r6.t0.t1.s4.clk ;
    wire [7:0] \AES.r6.t0.t1.s4.in ;
    reg [7:0] \AES.r6.t0.t1.s4.out ;
    wire \AES.r6.t0.t2.clk ;
    wire [7:0] \AES.r6.t0.t2.in ;
    wire [31:0] \AES.r6.t0.t2.out ;
    wire [7:0] \AES.r6.t0.t2.k0 ;
    wire [7:0] \AES.r6.t0.t2.k1 ;
    wire \AES.r6.t0.t2.s0.clk ;
    wire [7:0] \AES.r6.t0.t2.s0.in ;
    reg [7:0] \AES.r6.t0.t2.s0.out ;
    wire \AES.r6.t0.t2.s4.clk ;
    wire [7:0] \AES.r6.t0.t2.s4.in ;
    reg [7:0] \AES.r6.t0.t2.s4.out ;
    wire \AES.r6.t0.t3.clk ;
    wire [7:0] \AES.r6.t0.t3.in ;
    wire [31:0] \AES.r6.t0.t3.out ;
    wire [7:0] \AES.r6.t0.t3.k0 ;
    wire [7:0] \AES.r6.t0.t3.k1 ;
    wire \AES.r6.t0.t3.s0.clk ;
    wire [7:0] \AES.r6.t0.t3.s0.in ;
    reg [7:0] \AES.r6.t0.t3.s0.out ;
    wire \AES.r6.t0.t3.s4.clk ;
    wire [7:0] \AES.r6.t0.t3.s4.in ;
    reg [7:0] \AES.r6.t0.t3.s4.out ;
    wire \AES.r6.t1.clk ;
    wire [31:0] \AES.r6.t1.state ;
    wire [31:0] \AES.r6.t1.p0 ;
    wire [31:0] \AES.r6.t1.p1 ;
    wire [31:0] \AES.r6.t1.p2 ;
    wire [31:0] \AES.r6.t1.p3 ;
    wire [7:0] \AES.r6.t1.b0 ;
    wire [7:0] \AES.r6.t1.b1 ;
    wire [7:0] \AES.r6.t1.b2 ;
    wire [7:0] \AES.r6.t1.b3 ;
    wire [31:0] \AES.r6.t1.k0 ;
    wire [31:0] \AES.r6.t1.k1 ;
    wire [31:0] \AES.r6.t1.k2 ;
    wire \AES.r6.t1.t0.clk ;
    wire [7:0] \AES.r6.t1.t0.in ;
    wire [31:0] \AES.r6.t1.t0.out ;
    wire [7:0] \AES.r6.t1.t0.k0 ;
    wire [7:0] \AES.r6.t1.t0.k1 ;
    wire \AES.r6.t1.t0.s0.clk ;
    wire [7:0] \AES.r6.t1.t0.s0.in ;
    reg [7:0] \AES.r6.t1.t0.s0.out ;
    wire \AES.r6.t1.t0.s4.clk ;
    wire [7:0] \AES.r6.t1.t0.s4.in ;
    reg [7:0] \AES.r6.t1.t0.s4.out ;
    wire \AES.r6.t1.t1.clk ;
    wire [7:0] \AES.r6.t1.t1.in ;
    wire [31:0] \AES.r6.t1.t1.out ;
    wire [7:0] \AES.r6.t1.t1.k0 ;
    wire [7:0] \AES.r6.t1.t1.k1 ;
    wire \AES.r6.t1.t1.s0.clk ;
    wire [7:0] \AES.r6.t1.t1.s0.in ;
    reg [7:0] \AES.r6.t1.t1.s0.out ;
    wire \AES.r6.t1.t1.s4.clk ;
    wire [7:0] \AES.r6.t1.t1.s4.in ;
    reg [7:0] \AES.r6.t1.t1.s4.out ;
    wire \AES.r6.t1.t2.clk ;
    wire [7:0] \AES.r6.t1.t2.in ;
    wire [31:0] \AES.r6.t1.t2.out ;
    wire [7:0] \AES.r6.t1.t2.k0 ;
    wire [7:0] \AES.r6.t1.t2.k1 ;
    wire \AES.r6.t1.t2.s0.clk ;
    wire [7:0] \AES.r6.t1.t2.s0.in ;
    reg [7:0] \AES.r6.t1.t2.s0.out ;
    wire \AES.r6.t1.t2.s4.clk ;
    wire [7:0] \AES.r6.t1.t2.s4.in ;
    reg [7:0] \AES.r6.t1.t2.s4.out ;
    wire \AES.r6.t1.t3.clk ;
    wire [7:0] \AES.r6.t1.t3.in ;
    wire [31:0] \AES.r6.t1.t3.out ;
    wire [7:0] \AES.r6.t1.t3.k0 ;
    wire [7:0] \AES.r6.t1.t3.k1 ;
    wire \AES.r6.t1.t3.s0.clk ;
    wire [7:0] \AES.r6.t1.t3.s0.in ;
    reg [7:0] \AES.r6.t1.t3.s0.out ;
    wire \AES.r6.t1.t3.s4.clk ;
    wire [7:0] \AES.r6.t1.t3.s4.in ;
    reg [7:0] \AES.r6.t1.t3.s4.out ;
    wire \AES.r6.t2.clk ;
    wire [31:0] \AES.r6.t2.state ;
    wire [31:0] \AES.r6.t2.p0 ;
    wire [31:0] \AES.r6.t2.p1 ;
    wire [31:0] \AES.r6.t2.p2 ;
    wire [31:0] \AES.r6.t2.p3 ;
    wire [7:0] \AES.r6.t2.b0 ;
    wire [7:0] \AES.r6.t2.b1 ;
    wire [7:0] \AES.r6.t2.b2 ;
    wire [7:0] \AES.r6.t2.b3 ;
    wire [31:0] \AES.r6.t2.k0 ;
    wire [31:0] \AES.r6.t2.k1 ;
    wire [31:0] \AES.r6.t2.k2 ;
    wire \AES.r6.t2.t0.clk ;
    wire [7:0] \AES.r6.t2.t0.in ;
    wire [31:0] \AES.r6.t2.t0.out ;
    wire [7:0] \AES.r6.t2.t0.k0 ;
    wire [7:0] \AES.r6.t2.t0.k1 ;
    wire \AES.r6.t2.t0.s0.clk ;
    wire [7:0] \AES.r6.t2.t0.s0.in ;
    reg [7:0] \AES.r6.t2.t0.s0.out ;
    wire \AES.r6.t2.t0.s4.clk ;
    wire [7:0] \AES.r6.t2.t0.s4.in ;
    reg [7:0] \AES.r6.t2.t0.s4.out ;
    wire \AES.r6.t2.t1.clk ;
    wire [7:0] \AES.r6.t2.t1.in ;
    wire [31:0] \AES.r6.t2.t1.out ;
    wire [7:0] \AES.r6.t2.t1.k0 ;
    wire [7:0] \AES.r6.t2.t1.k1 ;
    wire \AES.r6.t2.t1.s0.clk ;
    wire [7:0] \AES.r6.t2.t1.s0.in ;
    reg [7:0] \AES.r6.t2.t1.s0.out ;
    wire \AES.r6.t2.t1.s4.clk ;
    wire [7:0] \AES.r6.t2.t1.s4.in ;
    reg [7:0] \AES.r6.t2.t1.s4.out ;
    wire \AES.r6.t2.t2.clk ;
    wire [7:0] \AES.r6.t2.t2.in ;
    wire [31:0] \AES.r6.t2.t2.out ;
    wire [7:0] \AES.r6.t2.t2.k0 ;
    wire [7:0] \AES.r6.t2.t2.k1 ;
    wire \AES.r6.t2.t2.s0.clk ;
    wire [7:0] \AES.r6.t2.t2.s0.in ;
    reg [7:0] \AES.r6.t2.t2.s0.out ;
    wire \AES.r6.t2.t2.s4.clk ;
    wire [7:0] \AES.r6.t2.t2.s4.in ;
    reg [7:0] \AES.r6.t2.t2.s4.out ;
    wire \AES.r6.t2.t3.clk ;
    wire [7:0] \AES.r6.t2.t3.in ;
    wire [31:0] \AES.r6.t2.t3.out ;
    wire [7:0] \AES.r6.t2.t3.k0 ;
    wire [7:0] \AES.r6.t2.t3.k1 ;
    wire \AES.r6.t2.t3.s0.clk ;
    wire [7:0] \AES.r6.t2.t3.s0.in ;
    reg [7:0] \AES.r6.t2.t3.s0.out ;
    wire \AES.r6.t2.t3.s4.clk ;
    wire [7:0] \AES.r6.t2.t3.s4.in ;
    reg [7:0] \AES.r6.t2.t3.s4.out ;
    wire \AES.r6.t3.clk ;
    wire [31:0] \AES.r6.t3.state ;
    wire [31:0] \AES.r6.t3.p0 ;
    wire [31:0] \AES.r6.t3.p1 ;
    wire [31:0] \AES.r6.t3.p2 ;
    wire [31:0] \AES.r6.t3.p3 ;
    wire [7:0] \AES.r6.t3.b0 ;
    wire [7:0] \AES.r6.t3.b1 ;
    wire [7:0] \AES.r6.t3.b2 ;
    wire [7:0] \AES.r6.t3.b3 ;
    wire [31:0] \AES.r6.t3.k0 ;
    wire [31:0] \AES.r6.t3.k1 ;
    wire [31:0] \AES.r6.t3.k2 ;
    wire \AES.r6.t3.t0.clk ;
    wire [7:0] \AES.r6.t3.t0.in ;
    wire [31:0] \AES.r6.t3.t0.out ;
    wire [7:0] \AES.r6.t3.t0.k0 ;
    wire [7:0] \AES.r6.t3.t0.k1 ;
    wire \AES.r6.t3.t0.s0.clk ;
    wire [7:0] \AES.r6.t3.t0.s0.in ;
    reg [7:0] \AES.r6.t3.t0.s0.out ;
    wire \AES.r6.t3.t0.s4.clk ;
    wire [7:0] \AES.r6.t3.t0.s4.in ;
    reg [7:0] \AES.r6.t3.t0.s4.out ;
    wire \AES.r6.t3.t1.clk ;
    wire [7:0] \AES.r6.t3.t1.in ;
    wire [31:0] \AES.r6.t3.t1.out ;
    wire [7:0] \AES.r6.t3.t1.k0 ;
    wire [7:0] \AES.r6.t3.t1.k1 ;
    wire \AES.r6.t3.t1.s0.clk ;
    wire [7:0] \AES.r6.t3.t1.s0.in ;
    reg [7:0] \AES.r6.t3.t1.s0.out ;
    wire \AES.r6.t3.t1.s4.clk ;
    wire [7:0] \AES.r6.t3.t1.s4.in ;
    reg [7:0] \AES.r6.t3.t1.s4.out ;
    wire \AES.r6.t3.t2.clk ;
    wire [7:0] \AES.r6.t3.t2.in ;
    wire [31:0] \AES.r6.t3.t2.out ;
    wire [7:0] \AES.r6.t3.t2.k0 ;
    wire [7:0] \AES.r6.t3.t2.k1 ;
    wire \AES.r6.t3.t2.s0.clk ;
    wire [7:0] \AES.r6.t3.t2.s0.in ;
    reg [7:0] \AES.r6.t3.t2.s0.out ;
    wire \AES.r6.t3.t2.s4.clk ;
    wire [7:0] \AES.r6.t3.t2.s4.in ;
    reg [7:0] \AES.r6.t3.t2.s4.out ;
    wire \AES.r6.t3.t3.clk ;
    wire [7:0] \AES.r6.t3.t3.in ;
    wire [31:0] \AES.r6.t3.t3.out ;
    wire [7:0] \AES.r6.t3.t3.k0 ;
    wire [7:0] \AES.r6.t3.t3.k1 ;
    wire \AES.r6.t3.t3.s0.clk ;
    wire [7:0] \AES.r6.t3.t3.s0.in ;
    reg [7:0] \AES.r6.t3.t3.s0.out ;
    wire \AES.r6.t3.t3.s4.clk ;
    wire [7:0] \AES.r6.t3.t3.s4.in ;
    reg [7:0] \AES.r6.t3.t3.s4.out ;
    wire \AES.r7.clk ;
    wire [127:0] \AES.r7.state_in ;
    wire [127:0] \AES.r7.key ;
    reg [127:0] \AES.r7.state_out ;
    wire [31:0] \AES.r7.s0 ;
    wire [31:0] \AES.r7.s1 ;
    wire [31:0] \AES.r7.s2 ;
    wire [31:0] \AES.r7.s3 ;
    wire [31:0] \AES.r7.z0 ;
    wire [31:0] \AES.r7.z1 ;
    wire [31:0] \AES.r7.z2 ;
    wire [31:0] \AES.r7.z3 ;
    wire [31:0] \AES.r7.p00 ;
    wire [31:0] \AES.r7.p01 ;
    wire [31:0] \AES.r7.p02 ;
    wire [31:0] \AES.r7.p03 ;
    wire [31:0] \AES.r7.p10 ;
    wire [31:0] \AES.r7.p11 ;
    wire [31:0] \AES.r7.p12 ;
    wire [31:0] \AES.r7.p13 ;
    wire [31:0] \AES.r7.p20 ;
    wire [31:0] \AES.r7.p21 ;
    wire [31:0] \AES.r7.p22 ;
    wire [31:0] \AES.r7.p23 ;
    wire [31:0] \AES.r7.p30 ;
    wire [31:0] \AES.r7.p31 ;
    wire [31:0] \AES.r7.p32 ;
    wire [31:0] \AES.r7.p33 ;
    wire [31:0] \AES.r7.k0 ;
    wire [31:0] \AES.r7.k1 ;
    wire [31:0] \AES.r7.k2 ;
    wire [31:0] \AES.r7.k3 ;
    wire \AES.r7.t0.clk ;
    wire [31:0] \AES.r7.t0.state ;
    wire [31:0] \AES.r7.t0.p0 ;
    wire [31:0] \AES.r7.t0.p1 ;
    wire [31:0] \AES.r7.t0.p2 ;
    wire [31:0] \AES.r7.t0.p3 ;
    wire [7:0] \AES.r7.t0.b0 ;
    wire [7:0] \AES.r7.t0.b1 ;
    wire [7:0] \AES.r7.t0.b2 ;
    wire [7:0] \AES.r7.t0.b3 ;
    wire [31:0] \AES.r7.t0.k0 ;
    wire [31:0] \AES.r7.t0.k1 ;
    wire [31:0] \AES.r7.t0.k2 ;
    wire \AES.r7.t0.t0.clk ;
    wire [7:0] \AES.r7.t0.t0.in ;
    wire [31:0] \AES.r7.t0.t0.out ;
    wire [7:0] \AES.r7.t0.t0.k0 ;
    wire [7:0] \AES.r7.t0.t0.k1 ;
    wire \AES.r7.t0.t0.s0.clk ;
    wire [7:0] \AES.r7.t0.t0.s0.in ;
    reg [7:0] \AES.r7.t0.t0.s0.out ;
    wire \AES.r7.t0.t0.s4.clk ;
    wire [7:0] \AES.r7.t0.t0.s4.in ;
    reg [7:0] \AES.r7.t0.t0.s4.out ;
    wire \AES.r7.t0.t1.clk ;
    wire [7:0] \AES.r7.t0.t1.in ;
    wire [31:0] \AES.r7.t0.t1.out ;
    wire [7:0] \AES.r7.t0.t1.k0 ;
    wire [7:0] \AES.r7.t0.t1.k1 ;
    wire \AES.r7.t0.t1.s0.clk ;
    wire [7:0] \AES.r7.t0.t1.s0.in ;
    reg [7:0] \AES.r7.t0.t1.s0.out ;
    wire \AES.r7.t0.t1.s4.clk ;
    wire [7:0] \AES.r7.t0.t1.s4.in ;
    reg [7:0] \AES.r7.t0.t1.s4.out ;
    wire \AES.r7.t0.t2.clk ;
    wire [7:0] \AES.r7.t0.t2.in ;
    wire [31:0] \AES.r7.t0.t2.out ;
    wire [7:0] \AES.r7.t0.t2.k0 ;
    wire [7:0] \AES.r7.t0.t2.k1 ;
    wire \AES.r7.t0.t2.s0.clk ;
    wire [7:0] \AES.r7.t0.t2.s0.in ;
    reg [7:0] \AES.r7.t0.t2.s0.out ;
    wire \AES.r7.t0.t2.s4.clk ;
    wire [7:0] \AES.r7.t0.t2.s4.in ;
    reg [7:0] \AES.r7.t0.t2.s4.out ;
    wire \AES.r7.t0.t3.clk ;
    wire [7:0] \AES.r7.t0.t3.in ;
    wire [31:0] \AES.r7.t0.t3.out ;
    wire [7:0] \AES.r7.t0.t3.k0 ;
    wire [7:0] \AES.r7.t0.t3.k1 ;
    wire \AES.r7.t0.t3.s0.clk ;
    wire [7:0] \AES.r7.t0.t3.s0.in ;
    reg [7:0] \AES.r7.t0.t3.s0.out ;
    wire \AES.r7.t0.t3.s4.clk ;
    wire [7:0] \AES.r7.t0.t3.s4.in ;
    reg [7:0] \AES.r7.t0.t3.s4.out ;
    wire \AES.r7.t1.clk ;
    wire [31:0] \AES.r7.t1.state ;
    wire [31:0] \AES.r7.t1.p0 ;
    wire [31:0] \AES.r7.t1.p1 ;
    wire [31:0] \AES.r7.t1.p2 ;
    wire [31:0] \AES.r7.t1.p3 ;
    wire [7:0] \AES.r7.t1.b0 ;
    wire [7:0] \AES.r7.t1.b1 ;
    wire [7:0] \AES.r7.t1.b2 ;
    wire [7:0] \AES.r7.t1.b3 ;
    wire [31:0] \AES.r7.t1.k0 ;
    wire [31:0] \AES.r7.t1.k1 ;
    wire [31:0] \AES.r7.t1.k2 ;
    wire \AES.r7.t1.t0.clk ;
    wire [7:0] \AES.r7.t1.t0.in ;
    wire [31:0] \AES.r7.t1.t0.out ;
    wire [7:0] \AES.r7.t1.t0.k0 ;
    wire [7:0] \AES.r7.t1.t0.k1 ;
    wire \AES.r7.t1.t0.s0.clk ;
    wire [7:0] \AES.r7.t1.t0.s0.in ;
    reg [7:0] \AES.r7.t1.t0.s0.out ;
    wire \AES.r7.t1.t0.s4.clk ;
    wire [7:0] \AES.r7.t1.t0.s4.in ;
    reg [7:0] \AES.r7.t1.t0.s4.out ;
    wire \AES.r7.t1.t1.clk ;
    wire [7:0] \AES.r7.t1.t1.in ;
    wire [31:0] \AES.r7.t1.t1.out ;
    wire [7:0] \AES.r7.t1.t1.k0 ;
    wire [7:0] \AES.r7.t1.t1.k1 ;
    wire \AES.r7.t1.t1.s0.clk ;
    wire [7:0] \AES.r7.t1.t1.s0.in ;
    reg [7:0] \AES.r7.t1.t1.s0.out ;
    wire \AES.r7.t1.t1.s4.clk ;
    wire [7:0] \AES.r7.t1.t1.s4.in ;
    reg [7:0] \AES.r7.t1.t1.s4.out ;
    wire \AES.r7.t1.t2.clk ;
    wire [7:0] \AES.r7.t1.t2.in ;
    wire [31:0] \AES.r7.t1.t2.out ;
    wire [7:0] \AES.r7.t1.t2.k0 ;
    wire [7:0] \AES.r7.t1.t2.k1 ;
    wire \AES.r7.t1.t2.s0.clk ;
    wire [7:0] \AES.r7.t1.t2.s0.in ;
    reg [7:0] \AES.r7.t1.t2.s0.out ;
    wire \AES.r7.t1.t2.s4.clk ;
    wire [7:0] \AES.r7.t1.t2.s4.in ;
    reg [7:0] \AES.r7.t1.t2.s4.out ;
    wire \AES.r7.t1.t3.clk ;
    wire [7:0] \AES.r7.t1.t3.in ;
    wire [31:0] \AES.r7.t1.t3.out ;
    wire [7:0] \AES.r7.t1.t3.k0 ;
    wire [7:0] \AES.r7.t1.t3.k1 ;
    wire \AES.r7.t1.t3.s0.clk ;
    wire [7:0] \AES.r7.t1.t3.s0.in ;
    reg [7:0] \AES.r7.t1.t3.s0.out ;
    wire \AES.r7.t1.t3.s4.clk ;
    wire [7:0] \AES.r7.t1.t3.s4.in ;
    reg [7:0] \AES.r7.t1.t3.s4.out ;
    wire \AES.r7.t2.clk ;
    wire [31:0] \AES.r7.t2.state ;
    wire [31:0] \AES.r7.t2.p0 ;
    wire [31:0] \AES.r7.t2.p1 ;
    wire [31:0] \AES.r7.t2.p2 ;
    wire [31:0] \AES.r7.t2.p3 ;
    wire [7:0] \AES.r7.t2.b0 ;
    wire [7:0] \AES.r7.t2.b1 ;
    wire [7:0] \AES.r7.t2.b2 ;
    wire [7:0] \AES.r7.t2.b3 ;
    wire [31:0] \AES.r7.t2.k0 ;
    wire [31:0] \AES.r7.t2.k1 ;
    wire [31:0] \AES.r7.t2.k2 ;
    wire \AES.r7.t2.t0.clk ;
    wire [7:0] \AES.r7.t2.t0.in ;
    wire [31:0] \AES.r7.t2.t0.out ;
    wire [7:0] \AES.r7.t2.t0.k0 ;
    wire [7:0] \AES.r7.t2.t0.k1 ;
    wire \AES.r7.t2.t0.s0.clk ;
    wire [7:0] \AES.r7.t2.t0.s0.in ;
    reg [7:0] \AES.r7.t2.t0.s0.out ;
    wire \AES.r7.t2.t0.s4.clk ;
    wire [7:0] \AES.r7.t2.t0.s4.in ;
    reg [7:0] \AES.r7.t2.t0.s4.out ;
    wire \AES.r7.t2.t1.clk ;
    wire [7:0] \AES.r7.t2.t1.in ;
    wire [31:0] \AES.r7.t2.t1.out ;
    wire [7:0] \AES.r7.t2.t1.k0 ;
    wire [7:0] \AES.r7.t2.t1.k1 ;
    wire \AES.r7.t2.t1.s0.clk ;
    wire [7:0] \AES.r7.t2.t1.s0.in ;
    reg [7:0] \AES.r7.t2.t1.s0.out ;
    wire \AES.r7.t2.t1.s4.clk ;
    wire [7:0] \AES.r7.t2.t1.s4.in ;
    reg [7:0] \AES.r7.t2.t1.s4.out ;
    wire \AES.r7.t2.t2.clk ;
    wire [7:0] \AES.r7.t2.t2.in ;
    wire [31:0] \AES.r7.t2.t2.out ;
    wire [7:0] \AES.r7.t2.t2.k0 ;
    wire [7:0] \AES.r7.t2.t2.k1 ;
    wire \AES.r7.t2.t2.s0.clk ;
    wire [7:0] \AES.r7.t2.t2.s0.in ;
    reg [7:0] \AES.r7.t2.t2.s0.out ;
    wire \AES.r7.t2.t2.s4.clk ;
    wire [7:0] \AES.r7.t2.t2.s4.in ;
    reg [7:0] \AES.r7.t2.t2.s4.out ;
    wire \AES.r7.t2.t3.clk ;
    wire [7:0] \AES.r7.t2.t3.in ;
    wire [31:0] \AES.r7.t2.t3.out ;
    wire [7:0] \AES.r7.t2.t3.k0 ;
    wire [7:0] \AES.r7.t2.t3.k1 ;
    wire \AES.r7.t2.t3.s0.clk ;
    wire [7:0] \AES.r7.t2.t3.s0.in ;
    reg [7:0] \AES.r7.t2.t3.s0.out ;
    wire \AES.r7.t2.t3.s4.clk ;
    wire [7:0] \AES.r7.t2.t3.s4.in ;
    reg [7:0] \AES.r7.t2.t3.s4.out ;
    wire \AES.r7.t3.clk ;
    wire [31:0] \AES.r7.t3.state ;
    wire [31:0] \AES.r7.t3.p0 ;
    wire [31:0] \AES.r7.t3.p1 ;
    wire [31:0] \AES.r7.t3.p2 ;
    wire [31:0] \AES.r7.t3.p3 ;
    wire [7:0] \AES.r7.t3.b0 ;
    wire [7:0] \AES.r7.t3.b1 ;
    wire [7:0] \AES.r7.t3.b2 ;
    wire [7:0] \AES.r7.t3.b3 ;
    wire [31:0] \AES.r7.t3.k0 ;
    wire [31:0] \AES.r7.t3.k1 ;
    wire [31:0] \AES.r7.t3.k2 ;
    wire \AES.r7.t3.t0.clk ;
    wire [7:0] \AES.r7.t3.t0.in ;
    wire [31:0] \AES.r7.t3.t0.out ;
    wire [7:0] \AES.r7.t3.t0.k0 ;
    wire [7:0] \AES.r7.t3.t0.k1 ;
    wire \AES.r7.t3.t0.s0.clk ;
    wire [7:0] \AES.r7.t3.t0.s0.in ;
    reg [7:0] \AES.r7.t3.t0.s0.out ;
    wire \AES.r7.t3.t0.s4.clk ;
    wire [7:0] \AES.r7.t3.t0.s4.in ;
    reg [7:0] \AES.r7.t3.t0.s4.out ;
    wire \AES.r7.t3.t1.clk ;
    wire [7:0] \AES.r7.t3.t1.in ;
    wire [31:0] \AES.r7.t3.t1.out ;
    wire [7:0] \AES.r7.t3.t1.k0 ;
    wire [7:0] \AES.r7.t3.t1.k1 ;
    wire \AES.r7.t3.t1.s0.clk ;
    wire [7:0] \AES.r7.t3.t1.s0.in ;
    reg [7:0] \AES.r7.t3.t1.s0.out ;
    wire \AES.r7.t3.t1.s4.clk ;
    wire [7:0] \AES.r7.t3.t1.s4.in ;
    reg [7:0] \AES.r7.t3.t1.s4.out ;
    wire \AES.r7.t3.t2.clk ;
    wire [7:0] \AES.r7.t3.t2.in ;
    wire [31:0] \AES.r7.t3.t2.out ;
    wire [7:0] \AES.r7.t3.t2.k0 ;
    wire [7:0] \AES.r7.t3.t2.k1 ;
    wire \AES.r7.t3.t2.s0.clk ;
    wire [7:0] \AES.r7.t3.t2.s0.in ;
    reg [7:0] \AES.r7.t3.t2.s0.out ;
    wire \AES.r7.t3.t2.s4.clk ;
    wire [7:0] \AES.r7.t3.t2.s4.in ;
    reg [7:0] \AES.r7.t3.t2.s4.out ;
    wire \AES.r7.t3.t3.clk ;
    wire [7:0] \AES.r7.t3.t3.in ;
    wire [31:0] \AES.r7.t3.t3.out ;
    wire [7:0] \AES.r7.t3.t3.k0 ;
    wire [7:0] \AES.r7.t3.t3.k1 ;
    wire \AES.r7.t3.t3.s0.clk ;
    wire [7:0] \AES.r7.t3.t3.s0.in ;
    reg [7:0] \AES.r7.t3.t3.s0.out ;
    wire \AES.r7.t3.t3.s4.clk ;
    wire [7:0] \AES.r7.t3.t3.s4.in ;
    reg [7:0] \AES.r7.t3.t3.s4.out ;
    wire \AES.r8.clk ;
    wire [127:0] \AES.r8.state_in ;
    wire [127:0] \AES.r8.key ;
    reg [127:0] \AES.r8.state_out ;
    wire [31:0] \AES.r8.s0 ;
    wire [31:0] \AES.r8.s1 ;
    wire [31:0] \AES.r8.s2 ;
    wire [31:0] \AES.r8.s3 ;
    wire [31:0] \AES.r8.z0 ;
    wire [31:0] \AES.r8.z1 ;
    wire [31:0] \AES.r8.z2 ;
    wire [31:0] \AES.r8.z3 ;
    wire [31:0] \AES.r8.p00 ;
    wire [31:0] \AES.r8.p01 ;
    wire [31:0] \AES.r8.p02 ;
    wire [31:0] \AES.r8.p03 ;
    wire [31:0] \AES.r8.p10 ;
    wire [31:0] \AES.r8.p11 ;
    wire [31:0] \AES.r8.p12 ;
    wire [31:0] \AES.r8.p13 ;
    wire [31:0] \AES.r8.p20 ;
    wire [31:0] \AES.r8.p21 ;
    wire [31:0] \AES.r8.p22 ;
    wire [31:0] \AES.r8.p23 ;
    wire [31:0] \AES.r8.p30 ;
    wire [31:0] \AES.r8.p31 ;
    wire [31:0] \AES.r8.p32 ;
    wire [31:0] \AES.r8.p33 ;
    wire [31:0] \AES.r8.k0 ;
    wire [31:0] \AES.r8.k1 ;
    wire [31:0] \AES.r8.k2 ;
    wire [31:0] \AES.r8.k3 ;
    wire \AES.r8.t0.clk ;
    wire [31:0] \AES.r8.t0.state ;
    wire [31:0] \AES.r8.t0.p0 ;
    wire [31:0] \AES.r8.t0.p1 ;
    wire [31:0] \AES.r8.t0.p2 ;
    wire [31:0] \AES.r8.t0.p3 ;
    wire [7:0] \AES.r8.t0.b0 ;
    wire [7:0] \AES.r8.t0.b1 ;
    wire [7:0] \AES.r8.t0.b2 ;
    wire [7:0] \AES.r8.t0.b3 ;
    wire [31:0] \AES.r8.t0.k0 ;
    wire [31:0] \AES.r8.t0.k1 ;
    wire [31:0] \AES.r8.t0.k2 ;
    wire \AES.r8.t0.t0.clk ;
    wire [7:0] \AES.r8.t0.t0.in ;
    wire [31:0] \AES.r8.t0.t0.out ;
    wire [7:0] \AES.r8.t0.t0.k0 ;
    wire [7:0] \AES.r8.t0.t0.k1 ;
    wire \AES.r8.t0.t0.s0.clk ;
    wire [7:0] \AES.r8.t0.t0.s0.in ;
    reg [7:0] \AES.r8.t0.t0.s0.out ;
    wire \AES.r8.t0.t0.s4.clk ;
    wire [7:0] \AES.r8.t0.t0.s4.in ;
    reg [7:0] \AES.r8.t0.t0.s4.out ;
    wire \AES.r8.t0.t1.clk ;
    wire [7:0] \AES.r8.t0.t1.in ;
    wire [31:0] \AES.r8.t0.t1.out ;
    wire [7:0] \AES.r8.t0.t1.k0 ;
    wire [7:0] \AES.r8.t0.t1.k1 ;
    wire \AES.r8.t0.t1.s0.clk ;
    wire [7:0] \AES.r8.t0.t1.s0.in ;
    reg [7:0] \AES.r8.t0.t1.s0.out ;
    wire \AES.r8.t0.t1.s4.clk ;
    wire [7:0] \AES.r8.t0.t1.s4.in ;
    reg [7:0] \AES.r8.t0.t1.s4.out ;
    wire \AES.r8.t0.t2.clk ;
    wire [7:0] \AES.r8.t0.t2.in ;
    wire [31:0] \AES.r8.t0.t2.out ;
    wire [7:0] \AES.r8.t0.t2.k0 ;
    wire [7:0] \AES.r8.t0.t2.k1 ;
    wire \AES.r8.t0.t2.s0.clk ;
    wire [7:0] \AES.r8.t0.t2.s0.in ;
    reg [7:0] \AES.r8.t0.t2.s0.out ;
    wire \AES.r8.t0.t2.s4.clk ;
    wire [7:0] \AES.r8.t0.t2.s4.in ;
    reg [7:0] \AES.r8.t0.t2.s4.out ;
    wire \AES.r8.t0.t3.clk ;
    wire [7:0] \AES.r8.t0.t3.in ;
    wire [31:0] \AES.r8.t0.t3.out ;
    wire [7:0] \AES.r8.t0.t3.k0 ;
    wire [7:0] \AES.r8.t0.t3.k1 ;
    wire \AES.r8.t0.t3.s0.clk ;
    wire [7:0] \AES.r8.t0.t3.s0.in ;
    reg [7:0] \AES.r8.t0.t3.s0.out ;
    wire \AES.r8.t0.t3.s4.clk ;
    wire [7:0] \AES.r8.t0.t3.s4.in ;
    reg [7:0] \AES.r8.t0.t3.s4.out ;
    wire \AES.r8.t1.clk ;
    wire [31:0] \AES.r8.t1.state ;
    wire [31:0] \AES.r8.t1.p0 ;
    wire [31:0] \AES.r8.t1.p1 ;
    wire [31:0] \AES.r8.t1.p2 ;
    wire [31:0] \AES.r8.t1.p3 ;
    wire [7:0] \AES.r8.t1.b0 ;
    wire [7:0] \AES.r8.t1.b1 ;
    wire [7:0] \AES.r8.t1.b2 ;
    wire [7:0] \AES.r8.t1.b3 ;
    wire [31:0] \AES.r8.t1.k0 ;
    wire [31:0] \AES.r8.t1.k1 ;
    wire [31:0] \AES.r8.t1.k2 ;
    wire \AES.r8.t1.t0.clk ;
    wire [7:0] \AES.r8.t1.t0.in ;
    wire [31:0] \AES.r8.t1.t0.out ;
    wire [7:0] \AES.r8.t1.t0.k0 ;
    wire [7:0] \AES.r8.t1.t0.k1 ;
    wire \AES.r8.t1.t0.s0.clk ;
    wire [7:0] \AES.r8.t1.t0.s0.in ;
    reg [7:0] \AES.r8.t1.t0.s0.out ;
    wire \AES.r8.t1.t0.s4.clk ;
    wire [7:0] \AES.r8.t1.t0.s4.in ;
    reg [7:0] \AES.r8.t1.t0.s4.out ;
    wire \AES.r8.t1.t1.clk ;
    wire [7:0] \AES.r8.t1.t1.in ;
    wire [31:0] \AES.r8.t1.t1.out ;
    wire [7:0] \AES.r8.t1.t1.k0 ;
    wire [7:0] \AES.r8.t1.t1.k1 ;
    wire \AES.r8.t1.t1.s0.clk ;
    wire [7:0] \AES.r8.t1.t1.s0.in ;
    reg [7:0] \AES.r8.t1.t1.s0.out ;
    wire \AES.r8.t1.t1.s4.clk ;
    wire [7:0] \AES.r8.t1.t1.s4.in ;
    reg [7:0] \AES.r8.t1.t1.s4.out ;
    wire \AES.r8.t1.t2.clk ;
    wire [7:0] \AES.r8.t1.t2.in ;
    wire [31:0] \AES.r8.t1.t2.out ;
    wire [7:0] \AES.r8.t1.t2.k0 ;
    wire [7:0] \AES.r8.t1.t2.k1 ;
    wire \AES.r8.t1.t2.s0.clk ;
    wire [7:0] \AES.r8.t1.t2.s0.in ;
    reg [7:0] \AES.r8.t1.t2.s0.out ;
    wire \AES.r8.t1.t2.s4.clk ;
    wire [7:0] \AES.r8.t1.t2.s4.in ;
    reg [7:0] \AES.r8.t1.t2.s4.out ;
    wire \AES.r8.t1.t3.clk ;
    wire [7:0] \AES.r8.t1.t3.in ;
    wire [31:0] \AES.r8.t1.t3.out ;
    wire [7:0] \AES.r8.t1.t3.k0 ;
    wire [7:0] \AES.r8.t1.t3.k1 ;
    wire \AES.r8.t1.t3.s0.clk ;
    wire [7:0] \AES.r8.t1.t3.s0.in ;
    reg [7:0] \AES.r8.t1.t3.s0.out ;
    wire \AES.r8.t1.t3.s4.clk ;
    wire [7:0] \AES.r8.t1.t3.s4.in ;
    reg [7:0] \AES.r8.t1.t3.s4.out ;
    wire \AES.r8.t2.clk ;
    wire [31:0] \AES.r8.t2.state ;
    wire [31:0] \AES.r8.t2.p0 ;
    wire [31:0] \AES.r8.t2.p1 ;
    wire [31:0] \AES.r8.t2.p2 ;
    wire [31:0] \AES.r8.t2.p3 ;
    wire [7:0] \AES.r8.t2.b0 ;
    wire [7:0] \AES.r8.t2.b1 ;
    wire [7:0] \AES.r8.t2.b2 ;
    wire [7:0] \AES.r8.t2.b3 ;
    wire [31:0] \AES.r8.t2.k0 ;
    wire [31:0] \AES.r8.t2.k1 ;
    wire [31:0] \AES.r8.t2.k2 ;
    wire \AES.r8.t2.t0.clk ;
    wire [7:0] \AES.r8.t2.t0.in ;
    wire [31:0] \AES.r8.t2.t0.out ;
    wire [7:0] \AES.r8.t2.t0.k0 ;
    wire [7:0] \AES.r8.t2.t0.k1 ;
    wire \AES.r8.t2.t0.s0.clk ;
    wire [7:0] \AES.r8.t2.t0.s0.in ;
    reg [7:0] \AES.r8.t2.t0.s0.out ;
    wire \AES.r8.t2.t0.s4.clk ;
    wire [7:0] \AES.r8.t2.t0.s4.in ;
    reg [7:0] \AES.r8.t2.t0.s4.out ;
    wire \AES.r8.t2.t1.clk ;
    wire [7:0] \AES.r8.t2.t1.in ;
    wire [31:0] \AES.r8.t2.t1.out ;
    wire [7:0] \AES.r8.t2.t1.k0 ;
    wire [7:0] \AES.r8.t2.t1.k1 ;
    wire \AES.r8.t2.t1.s0.clk ;
    wire [7:0] \AES.r8.t2.t1.s0.in ;
    reg [7:0] \AES.r8.t2.t1.s0.out ;
    wire \AES.r8.t2.t1.s4.clk ;
    wire [7:0] \AES.r8.t2.t1.s4.in ;
    reg [7:0] \AES.r8.t2.t1.s4.out ;
    wire \AES.r8.t2.t2.clk ;
    wire [7:0] \AES.r8.t2.t2.in ;
    wire [31:0] \AES.r8.t2.t2.out ;
    wire [7:0] \AES.r8.t2.t2.k0 ;
    wire [7:0] \AES.r8.t2.t2.k1 ;
    wire \AES.r8.t2.t2.s0.clk ;
    wire [7:0] \AES.r8.t2.t2.s0.in ;
    reg [7:0] \AES.r8.t2.t2.s0.out ;
    wire \AES.r8.t2.t2.s4.clk ;
    wire [7:0] \AES.r8.t2.t2.s4.in ;
    reg [7:0] \AES.r8.t2.t2.s4.out ;
    wire \AES.r8.t2.t3.clk ;
    wire [7:0] \AES.r8.t2.t3.in ;
    wire [31:0] \AES.r8.t2.t3.out ;
    wire [7:0] \AES.r8.t2.t3.k0 ;
    wire [7:0] \AES.r8.t2.t3.k1 ;
    wire \AES.r8.t2.t3.s0.clk ;
    wire [7:0] \AES.r8.t2.t3.s0.in ;
    reg [7:0] \AES.r8.t2.t3.s0.out ;
    wire \AES.r8.t2.t3.s4.clk ;
    wire [7:0] \AES.r8.t2.t3.s4.in ;
    reg [7:0] \AES.r8.t2.t3.s4.out ;
    wire \AES.r8.t3.clk ;
    wire [31:0] \AES.r8.t3.state ;
    wire [31:0] \AES.r8.t3.p0 ;
    wire [31:0] \AES.r8.t3.p1 ;
    wire [31:0] \AES.r8.t3.p2 ;
    wire [31:0] \AES.r8.t3.p3 ;
    wire [7:0] \AES.r8.t3.b0 ;
    wire [7:0] \AES.r8.t3.b1 ;
    wire [7:0] \AES.r8.t3.b2 ;
    wire [7:0] \AES.r8.t3.b3 ;
    wire [31:0] \AES.r8.t3.k0 ;
    wire [31:0] \AES.r8.t3.k1 ;
    wire [31:0] \AES.r8.t3.k2 ;
    wire \AES.r8.t3.t0.clk ;
    wire [7:0] \AES.r8.t3.t0.in ;
    wire [31:0] \AES.r8.t3.t0.out ;
    wire [7:0] \AES.r8.t3.t0.k0 ;
    wire [7:0] \AES.r8.t3.t0.k1 ;
    wire \AES.r8.t3.t0.s0.clk ;
    wire [7:0] \AES.r8.t3.t0.s0.in ;
    reg [7:0] \AES.r8.t3.t0.s0.out ;
    wire \AES.r8.t3.t0.s4.clk ;
    wire [7:0] \AES.r8.t3.t0.s4.in ;
    reg [7:0] \AES.r8.t3.t0.s4.out ;
    wire \AES.r8.t3.t1.clk ;
    wire [7:0] \AES.r8.t3.t1.in ;
    wire [31:0] \AES.r8.t3.t1.out ;
    wire [7:0] \AES.r8.t3.t1.k0 ;
    wire [7:0] \AES.r8.t3.t1.k1 ;
    wire \AES.r8.t3.t1.s0.clk ;
    wire [7:0] \AES.r8.t3.t1.s0.in ;
    reg [7:0] \AES.r8.t3.t1.s0.out ;
    wire \AES.r8.t3.t1.s4.clk ;
    wire [7:0] \AES.r8.t3.t1.s4.in ;
    reg [7:0] \AES.r8.t3.t1.s4.out ;
    wire \AES.r8.t3.t2.clk ;
    wire [7:0] \AES.r8.t3.t2.in ;
    wire [31:0] \AES.r8.t3.t2.out ;
    wire [7:0] \AES.r8.t3.t2.k0 ;
    wire [7:0] \AES.r8.t3.t2.k1 ;
    wire \AES.r8.t3.t2.s0.clk ;
    wire [7:0] \AES.r8.t3.t2.s0.in ;
    reg [7:0] \AES.r8.t3.t2.s0.out ;
    wire \AES.r8.t3.t2.s4.clk ;
    wire [7:0] \AES.r8.t3.t2.s4.in ;
    reg [7:0] \AES.r8.t3.t2.s4.out ;
    wire \AES.r8.t3.t3.clk ;
    wire [7:0] \AES.r8.t3.t3.in ;
    wire [31:0] \AES.r8.t3.t3.out ;
    wire [7:0] \AES.r8.t3.t3.k0 ;
    wire [7:0] \AES.r8.t3.t3.k1 ;
    wire \AES.r8.t3.t3.s0.clk ;
    wire [7:0] \AES.r8.t3.t3.s0.in ;
    reg [7:0] \AES.r8.t3.t3.s0.out ;
    wire \AES.r8.t3.t3.s4.clk ;
    wire [7:0] \AES.r8.t3.t3.s4.in ;
    reg [7:0] \AES.r8.t3.t3.s4.out ;
    wire \AES.r9.clk ;
    wire [127:0] \AES.r9.state_in ;
    wire [127:0] \AES.r9.key ;
    reg [127:0] \AES.r9.state_out ;
    wire [31:0] \AES.r9.s0 ;
    wire [31:0] \AES.r9.s1 ;
    wire [31:0] \AES.r9.s2 ;
    wire [31:0] \AES.r9.s3 ;
    wire [31:0] \AES.r9.z0 ;
    wire [31:0] \AES.r9.z1 ;
    wire [31:0] \AES.r9.z2 ;
    wire [31:0] \AES.r9.z3 ;
    wire [31:0] \AES.r9.p00 ;
    wire [31:0] \AES.r9.p01 ;
    wire [31:0] \AES.r9.p02 ;
    wire [31:0] \AES.r9.p03 ;
    wire [31:0] \AES.r9.p10 ;
    wire [31:0] \AES.r9.p11 ;
    wire [31:0] \AES.r9.p12 ;
    wire [31:0] \AES.r9.p13 ;
    wire [31:0] \AES.r9.p20 ;
    wire [31:0] \AES.r9.p21 ;
    wire [31:0] \AES.r9.p22 ;
    wire [31:0] \AES.r9.p23 ;
    wire [31:0] \AES.r9.p30 ;
    wire [31:0] \AES.r9.p31 ;
    wire [31:0] \AES.r9.p32 ;
    wire [31:0] \AES.r9.p33 ;
    wire [31:0] \AES.r9.k0 ;
    wire [31:0] \AES.r9.k1 ;
    wire [31:0] \AES.r9.k2 ;
    wire [31:0] \AES.r9.k3 ;
    wire \AES.r9.t0.clk ;
    wire [31:0] \AES.r9.t0.state ;
    wire [31:0] \AES.r9.t0.p0 ;
    wire [31:0] \AES.r9.t0.p1 ;
    wire [31:0] \AES.r9.t0.p2 ;
    wire [31:0] \AES.r9.t0.p3 ;
    wire [7:0] \AES.r9.t0.b0 ;
    wire [7:0] \AES.r9.t0.b1 ;
    wire [7:0] \AES.r9.t0.b2 ;
    wire [7:0] \AES.r9.t0.b3 ;
    wire [31:0] \AES.r9.t0.k0 ;
    wire [31:0] \AES.r9.t0.k1 ;
    wire [31:0] \AES.r9.t0.k2 ;
    wire \AES.r9.t0.t0.clk ;
    wire [7:0] \AES.r9.t0.t0.in ;
    wire [31:0] \AES.r9.t0.t0.out ;
    wire [7:0] \AES.r9.t0.t0.k0 ;
    wire [7:0] \AES.r9.t0.t0.k1 ;
    wire \AES.r9.t0.t0.s0.clk ;
    wire [7:0] \AES.r9.t0.t0.s0.in ;
    reg [7:0] \AES.r9.t0.t0.s0.out ;
    wire \AES.r9.t0.t0.s4.clk ;
    wire [7:0] \AES.r9.t0.t0.s4.in ;
    reg [7:0] \AES.r9.t0.t0.s4.out ;
    wire \AES.r9.t0.t1.clk ;
    wire [7:0] \AES.r9.t0.t1.in ;
    wire [31:0] \AES.r9.t0.t1.out ;
    wire [7:0] \AES.r9.t0.t1.k0 ;
    wire [7:0] \AES.r9.t0.t1.k1 ;
    wire \AES.r9.t0.t1.s0.clk ;
    wire [7:0] \AES.r9.t0.t1.s0.in ;
    reg [7:0] \AES.r9.t0.t1.s0.out ;
    wire \AES.r9.t0.t1.s4.clk ;
    wire [7:0] \AES.r9.t0.t1.s4.in ;
    reg [7:0] \AES.r9.t0.t1.s4.out ;
    wire \AES.r9.t0.t2.clk ;
    wire [7:0] \AES.r9.t0.t2.in ;
    wire [31:0] \AES.r9.t0.t2.out ;
    wire [7:0] \AES.r9.t0.t2.k0 ;
    wire [7:0] \AES.r9.t0.t2.k1 ;
    wire \AES.r9.t0.t2.s0.clk ;
    wire [7:0] \AES.r9.t0.t2.s0.in ;
    reg [7:0] \AES.r9.t0.t2.s0.out ;
    wire \AES.r9.t0.t2.s4.clk ;
    wire [7:0] \AES.r9.t0.t2.s4.in ;
    reg [7:0] \AES.r9.t0.t2.s4.out ;
    wire \AES.r9.t0.t3.clk ;
    wire [7:0] \AES.r9.t0.t3.in ;
    wire [31:0] \AES.r9.t0.t3.out ;
    wire [7:0] \AES.r9.t0.t3.k0 ;
    wire [7:0] \AES.r9.t0.t3.k1 ;
    wire \AES.r9.t0.t3.s0.clk ;
    wire [7:0] \AES.r9.t0.t3.s0.in ;
    reg [7:0] \AES.r9.t0.t3.s0.out ;
    wire \AES.r9.t0.t3.s4.clk ;
    wire [7:0] \AES.r9.t0.t3.s4.in ;
    reg [7:0] \AES.r9.t0.t3.s4.out ;
    wire \AES.r9.t1.clk ;
    wire [31:0] \AES.r9.t1.state ;
    wire [31:0] \AES.r9.t1.p0 ;
    wire [31:0] \AES.r9.t1.p1 ;
    wire [31:0] \AES.r9.t1.p2 ;
    wire [31:0] \AES.r9.t1.p3 ;
    wire [7:0] \AES.r9.t1.b0 ;
    wire [7:0] \AES.r9.t1.b1 ;
    wire [7:0] \AES.r9.t1.b2 ;
    wire [7:0] \AES.r9.t1.b3 ;
    wire [31:0] \AES.r9.t1.k0 ;
    wire [31:0] \AES.r9.t1.k1 ;
    wire [31:0] \AES.r9.t1.k2 ;
    wire \AES.r9.t1.t0.clk ;
    wire [7:0] \AES.r9.t1.t0.in ;
    wire [31:0] \AES.r9.t1.t0.out ;
    wire [7:0] \AES.r9.t1.t0.k0 ;
    wire [7:0] \AES.r9.t1.t0.k1 ;
    wire \AES.r9.t1.t0.s0.clk ;
    wire [7:0] \AES.r9.t1.t0.s0.in ;
    reg [7:0] \AES.r9.t1.t0.s0.out ;
    wire \AES.r9.t1.t0.s4.clk ;
    wire [7:0] \AES.r9.t1.t0.s4.in ;
    reg [7:0] \AES.r9.t1.t0.s4.out ;
    wire \AES.r9.t1.t1.clk ;
    wire [7:0] \AES.r9.t1.t1.in ;
    wire [31:0] \AES.r9.t1.t1.out ;
    wire [7:0] \AES.r9.t1.t1.k0 ;
    wire [7:0] \AES.r9.t1.t1.k1 ;
    wire \AES.r9.t1.t1.s0.clk ;
    wire [7:0] \AES.r9.t1.t1.s0.in ;
    reg [7:0] \AES.r9.t1.t1.s0.out ;
    wire \AES.r9.t1.t1.s4.clk ;
    wire [7:0] \AES.r9.t1.t1.s4.in ;
    reg [7:0] \AES.r9.t1.t1.s4.out ;
    wire \AES.r9.t1.t2.clk ;
    wire [7:0] \AES.r9.t1.t2.in ;
    wire [31:0] \AES.r9.t1.t2.out ;
    wire [7:0] \AES.r9.t1.t2.k0 ;
    wire [7:0] \AES.r9.t1.t2.k1 ;
    wire \AES.r9.t1.t2.s0.clk ;
    wire [7:0] \AES.r9.t1.t2.s0.in ;
    reg [7:0] \AES.r9.t1.t2.s0.out ;
    wire \AES.r9.t1.t2.s4.clk ;
    wire [7:0] \AES.r9.t1.t2.s4.in ;
    reg [7:0] \AES.r9.t1.t2.s4.out ;
    wire \AES.r9.t1.t3.clk ;
    wire [7:0] \AES.r9.t1.t3.in ;
    wire [31:0] \AES.r9.t1.t3.out ;
    wire [7:0] \AES.r9.t1.t3.k0 ;
    wire [7:0] \AES.r9.t1.t3.k1 ;
    wire \AES.r9.t1.t3.s0.clk ;
    wire [7:0] \AES.r9.t1.t3.s0.in ;
    reg [7:0] \AES.r9.t1.t3.s0.out ;
    wire \AES.r9.t1.t3.s4.clk ;
    wire [7:0] \AES.r9.t1.t3.s4.in ;
    reg [7:0] \AES.r9.t1.t3.s4.out ;
    wire \AES.r9.t2.clk ;
    wire [31:0] \AES.r9.t2.state ;
    wire [31:0] \AES.r9.t2.p0 ;
    wire [31:0] \AES.r9.t2.p1 ;
    wire [31:0] \AES.r9.t2.p2 ;
    wire [31:0] \AES.r9.t2.p3 ;
    wire [7:0] \AES.r9.t2.b0 ;
    wire [7:0] \AES.r9.t2.b1 ;
    wire [7:0] \AES.r9.t2.b2 ;
    wire [7:0] \AES.r9.t2.b3 ;
    wire [31:0] \AES.r9.t2.k0 ;
    wire [31:0] \AES.r9.t2.k1 ;
    wire [31:0] \AES.r9.t2.k2 ;
    wire \AES.r9.t2.t0.clk ;
    wire [7:0] \AES.r9.t2.t0.in ;
    wire [31:0] \AES.r9.t2.t0.out ;
    wire [7:0] \AES.r9.t2.t0.k0 ;
    wire [7:0] \AES.r9.t2.t0.k1 ;
    wire \AES.r9.t2.t0.s0.clk ;
    wire [7:0] \AES.r9.t2.t0.s0.in ;
    reg [7:0] \AES.r9.t2.t0.s0.out ;
    wire \AES.r9.t2.t0.s4.clk ;
    wire [7:0] \AES.r9.t2.t0.s4.in ;
    reg [7:0] \AES.r9.t2.t0.s4.out ;
    wire \AES.r9.t2.t1.clk ;
    wire [7:0] \AES.r9.t2.t1.in ;
    wire [31:0] \AES.r9.t2.t1.out ;
    wire [7:0] \AES.r9.t2.t1.k0 ;
    wire [7:0] \AES.r9.t2.t1.k1 ;
    wire \AES.r9.t2.t1.s0.clk ;
    wire [7:0] \AES.r9.t2.t1.s0.in ;
    reg [7:0] \AES.r9.t2.t1.s0.out ;
    wire \AES.r9.t2.t1.s4.clk ;
    wire [7:0] \AES.r9.t2.t1.s4.in ;
    reg [7:0] \AES.r9.t2.t1.s4.out ;
    wire \AES.r9.t2.t2.clk ;
    wire [7:0] \AES.r9.t2.t2.in ;
    wire [31:0] \AES.r9.t2.t2.out ;
    wire [7:0] \AES.r9.t2.t2.k0 ;
    wire [7:0] \AES.r9.t2.t2.k1 ;
    wire \AES.r9.t2.t2.s0.clk ;
    wire [7:0] \AES.r9.t2.t2.s0.in ;
    reg [7:0] \AES.r9.t2.t2.s0.out ;
    wire \AES.r9.t2.t2.s4.clk ;
    wire [7:0] \AES.r9.t2.t2.s4.in ;
    reg [7:0] \AES.r9.t2.t2.s4.out ;
    wire \AES.r9.t2.t3.clk ;
    wire [7:0] \AES.r9.t2.t3.in ;
    wire [31:0] \AES.r9.t2.t3.out ;
    wire [7:0] \AES.r9.t2.t3.k0 ;
    wire [7:0] \AES.r9.t2.t3.k1 ;
    wire \AES.r9.t2.t3.s0.clk ;
    wire [7:0] \AES.r9.t2.t3.s0.in ;
    reg [7:0] \AES.r9.t2.t3.s0.out ;
    wire \AES.r9.t2.t3.s4.clk ;
    wire [7:0] \AES.r9.t2.t3.s4.in ;
    reg [7:0] \AES.r9.t2.t3.s4.out ;
    wire \AES.r9.t3.clk ;
    wire [31:0] \AES.r9.t3.state ;
    wire [31:0] \AES.r9.t3.p0 ;
    wire [31:0] \AES.r9.t3.p1 ;
    wire [31:0] \AES.r9.t3.p2 ;
    wire [31:0] \AES.r9.t3.p3 ;
    wire [7:0] \AES.r9.t3.b0 ;
    wire [7:0] \AES.r9.t3.b1 ;
    wire [7:0] \AES.r9.t3.b2 ;
    wire [7:0] \AES.r9.t3.b3 ;
    wire [31:0] \AES.r9.t3.k0 ;
    wire [31:0] \AES.r9.t3.k1 ;
    wire [31:0] \AES.r9.t3.k2 ;
    wire \AES.r9.t3.t0.clk ;
    wire [7:0] \AES.r9.t3.t0.in ;
    wire [31:0] \AES.r9.t3.t0.out ;
    wire [7:0] \AES.r9.t3.t0.k0 ;
    wire [7:0] \AES.r9.t3.t0.k1 ;
    wire \AES.r9.t3.t0.s0.clk ;
    wire [7:0] \AES.r9.t3.t0.s0.in ;
    reg [7:0] \AES.r9.t3.t0.s0.out ;
    wire \AES.r9.t3.t0.s4.clk ;
    wire [7:0] \AES.r9.t3.t0.s4.in ;
    reg [7:0] \AES.r9.t3.t0.s4.out ;
    wire \AES.r9.t3.t1.clk ;
    wire [7:0] \AES.r9.t3.t1.in ;
    wire [31:0] \AES.r9.t3.t1.out ;
    wire [7:0] \AES.r9.t3.t1.k0 ;
    wire [7:0] \AES.r9.t3.t1.k1 ;
    wire \AES.r9.t3.t1.s0.clk ;
    wire [7:0] \AES.r9.t3.t1.s0.in ;
    reg [7:0] \AES.r9.t3.t1.s0.out ;
    wire \AES.r9.t3.t1.s4.clk ;
    wire [7:0] \AES.r9.t3.t1.s4.in ;
    reg [7:0] \AES.r9.t3.t1.s4.out ;
    wire \AES.r9.t3.t2.clk ;
    wire [7:0] \AES.r9.t3.t2.in ;
    wire [31:0] \AES.r9.t3.t2.out ;
    wire [7:0] \AES.r9.t3.t2.k0 ;
    wire [7:0] \AES.r9.t3.t2.k1 ;
    wire \AES.r9.t3.t2.s0.clk ;
    wire [7:0] \AES.r9.t3.t2.s0.in ;
    reg [7:0] \AES.r9.t3.t2.s0.out ;
    wire \AES.r9.t3.t2.s4.clk ;
    wire [7:0] \AES.r9.t3.t2.s4.in ;
    reg [7:0] \AES.r9.t3.t2.s4.out ;
    wire \AES.r9.t3.t3.clk ;
    wire [7:0] \AES.r9.t3.t3.in ;
    wire [31:0] \AES.r9.t3.t3.out ;
    wire [7:0] \AES.r9.t3.t3.k0 ;
    wire [7:0] \AES.r9.t3.t3.k1 ;
    wire \AES.r9.t3.t3.s0.clk ;
    wire [7:0] \AES.r9.t3.t3.s0.in ;
    reg [7:0] \AES.r9.t3.t3.s0.out ;
    wire \AES.r9.t3.t3.s4.clk ;
    wire [7:0] \AES.r9.t3.t3.s4.in ;
    reg [7:0] \AES.r9.t3.t3.s4.out ;
    wire \AES.rf.clk ;
    wire [127:0] \AES.rf.state_in ;
    wire [127:0] \AES.rf.key_in ;
    reg [127:0] \AES.rf.state_out ;
    wire [31:0] \AES.rf.s0 ;
    wire [31:0] \AES.rf.s1 ;
    wire [31:0] \AES.rf.s2 ;
    wire [31:0] \AES.rf.s3 ;
    wire [31:0] \AES.rf.z0 ;
    wire [31:0] \AES.rf.z1 ;
    wire [31:0] \AES.rf.z2 ;
    wire [31:0] \AES.rf.z3 ;
    wire [31:0] \AES.rf.k0 ;
    wire [31:0] \AES.rf.k1 ;
    wire [31:0] \AES.rf.k2 ;
    wire [31:0] \AES.rf.k3 ;
    wire [7:0] \AES.rf.p00 ;
    wire [7:0] \AES.rf.p01 ;
    wire [7:0] \AES.rf.p02 ;
    wire [7:0] \AES.rf.p03 ;
    wire [7:0] \AES.rf.p10 ;
    wire [7:0] \AES.rf.p11 ;
    wire [7:0] \AES.rf.p12 ;
    wire [7:0] \AES.rf.p13 ;
    wire [7:0] \AES.rf.p20 ;
    wire [7:0] \AES.rf.p21 ;
    wire [7:0] \AES.rf.p22 ;
    wire [7:0] \AES.rf.p23 ;
    wire [7:0] \AES.rf.p30 ;
    wire [7:0] \AES.rf.p31 ;
    wire [7:0] \AES.rf.p32 ;
    wire [7:0] \AES.rf.p33 ;
    wire \AES.rf.S4_1.clk ;
    wire [31:0] \AES.rf.S4_1.in ;
    wire [31:0] \AES.rf.S4_1.out ;
    wire [7:0] \AES.rf.S4_1.k0 ;
    wire [7:0] \AES.rf.S4_1.k1 ;
    wire [7:0] \AES.rf.S4_1.k2 ;
    wire [7:0] \AES.rf.S4_1.k3 ;
    wire \AES.rf.S4_1.S_0.clk ;
    wire [7:0] \AES.rf.S4_1.S_0.in ;
    reg [7:0] \AES.rf.S4_1.S_0.out ;
    wire \AES.rf.S4_1.S_1.clk ;
    wire [7:0] \AES.rf.S4_1.S_1.in ;
    reg [7:0] \AES.rf.S4_1.S_1.out ;
    wire \AES.rf.S4_1.S_2.clk ;
    wire [7:0] \AES.rf.S4_1.S_2.in ;
    reg [7:0] \AES.rf.S4_1.S_2.out ;
    wire \AES.rf.S4_1.S_3.clk ;
    wire [7:0] \AES.rf.S4_1.S_3.in ;
    reg [7:0] \AES.rf.S4_1.S_3.out ;
    wire \AES.rf.S4_2.clk ;
    wire [31:0] \AES.rf.S4_2.in ;
    wire [31:0] \AES.rf.S4_2.out ;
    wire [7:0] \AES.rf.S4_2.k0 ;
    wire [7:0] \AES.rf.S4_2.k1 ;
    wire [7:0] \AES.rf.S4_2.k2 ;
    wire [7:0] \AES.rf.S4_2.k3 ;
    wire \AES.rf.S4_2.S_0.clk ;
    wire [7:0] \AES.rf.S4_2.S_0.in ;
    reg [7:0] \AES.rf.S4_2.S_0.out ;
    wire \AES.rf.S4_2.S_1.clk ;
    wire [7:0] \AES.rf.S4_2.S_1.in ;
    reg [7:0] \AES.rf.S4_2.S_1.out ;
    wire \AES.rf.S4_2.S_2.clk ;
    wire [7:0] \AES.rf.S4_2.S_2.in ;
    reg [7:0] \AES.rf.S4_2.S_2.out ;
    wire \AES.rf.S4_2.S_3.clk ;
    wire [7:0] \AES.rf.S4_2.S_3.in ;
    reg [7:0] \AES.rf.S4_2.S_3.out ;
    wire \AES.rf.S4_3.clk ;
    wire [31:0] \AES.rf.S4_3.in ;
    wire [31:0] \AES.rf.S4_3.out ;
    wire [7:0] \AES.rf.S4_3.k0 ;
    wire [7:0] \AES.rf.S4_3.k1 ;
    wire [7:0] \AES.rf.S4_3.k2 ;
    wire [7:0] \AES.rf.S4_3.k3 ;
    wire \AES.rf.S4_3.S_0.clk ;
    wire [7:0] \AES.rf.S4_3.S_0.in ;
    reg [7:0] \AES.rf.S4_3.S_0.out ;
    wire \AES.rf.S4_3.S_1.clk ;
    wire [7:0] \AES.rf.S4_3.S_1.in ;
    reg [7:0] \AES.rf.S4_3.S_1.out ;
    wire \AES.rf.S4_3.S_2.clk ;
    wire [7:0] \AES.rf.S4_3.S_2.in ;
    reg [7:0] \AES.rf.S4_3.S_2.out ;
    wire \AES.rf.S4_3.S_3.clk ;
    wire [7:0] \AES.rf.S4_3.S_3.in ;
    reg [7:0] \AES.rf.S4_3.S_3.out ;
    wire \AES.rf.S4_4.clk ;
    wire [31:0] \AES.rf.S4_4.in ;
    wire [31:0] \AES.rf.S4_4.out ;
    wire [7:0] \AES.rf.S4_4.k0 ;
    wire [7:0] \AES.rf.S4_4.k1 ;
    wire [7:0] \AES.rf.S4_4.k2 ;
    wire [7:0] \AES.rf.S4_4.k3 ;
    wire \AES.rf.S4_4.S_0.clk ;
    wire [7:0] \AES.rf.S4_4.S_0.in ;
    reg [7:0] \AES.rf.S4_4.S_0.out ;
    wire \AES.rf.S4_4.S_1.clk ;
    wire [7:0] \AES.rf.S4_4.S_1.in ;
    reg [7:0] \AES.rf.S4_4.S_1.out ;
    wire \AES.rf.S4_4.S_2.clk ;
    wire [7:0] \AES.rf.S4_4.S_2.in ;
    reg [7:0] \AES.rf.S4_4.S_2.out ;
    wire \AES.rf.S4_4.S_3.clk ;
    wire [7:0] \AES.rf.S4_4.S_3.in ;
    reg [7:0] \AES.rf.S4_4.S_3.out ;
    assign \AES.clk  = clk;
    assign \AES.state  = state;
    assign \AES.key  = key;
    assign out = \AES.out ;
    always @ (  posedge \AES.clk )
    begin
        \AES.s0  <= ( \AES.state  ^ \AES.key  );
        \AES.k0  <= \AES.key ;
    end
    assign \AES.a1.clk  = \AES.clk ;
    assign \AES.a1.in  = \AES.k0 ;
    assign \AES.a1.rcon  = \AES.k1 ;
    assign \AES.k0b  = \AES.a1.out_1 ;
    assign \AES.a1_rcon  = \AES.a1.out_2 ;
    assign \AES.a1.k0  = \AES.a1.in [127:96];
    assign \AES.a1.k1  = \AES.a1.in [95:64];
    assign \AES.a1.k2  = \AES.a1.in [63:32];
    assign \AES.a1.k3  = \AES.a1.in [31:0];
    assign \AES.a1.v0  = { ( \AES.a1.k0 [31:24] ^ \AES.a1.rcon  ), \AES.a1.k0 [23:0] };
    assign \AES.a1.v1  = ( \AES.a1.v0  ^ \AES.a1.k1  );
    assign \AES.a1.v2  = ( \AES.a1.v1  ^ \AES.a1.k2  );
    assign \AES.a1.v3  = ( \AES.a1.v2  ^ \AES.a1.k3  );
    always @ (  posedge \AES.a1.clk )
    begin
        \AES.a1.k0a  <= \AES.a1.v0 ;
        \AES.a1.k1a  <= \AES.a1.v1 ;
        \AES.a1.k2a  <= \AES.a1.v2 ;
        \AES.a1.k3a  <= \AES.a1.v3 ;
    end
    assign \AES.a1.S4_0.clk  = \AES.a1.clk ;
    assign \AES.a1.S4_0.in  = { \AES.a1.k3 [23:0], \AES.a1.k3 [31:24] };
    assign \AES.a1.k4a  = \AES.a1.S4_0.out ;
    assign \AES.a1.S4_0.S_0.clk  = \AES.a1.S4_0.clk ;
    assign \AES.a1.S4_0.S_0.in  = \AES.a1.S4_0.in [31:24];
    assign \AES.a1.S4_0.k0  = \AES.a1.S4_0.S_0.out ;
    always @ (  posedge \AES.a1.S4_0.S_0.clk )
    begin
        case ( \AES.a1.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a1.S4_0.S_1.clk  = \AES.a1.S4_0.clk ;
    assign \AES.a1.S4_0.S_1.in  = \AES.a1.S4_0.in [23:16];
    assign \AES.a1.S4_0.k1  = \AES.a1.S4_0.S_1.out ;
    always @ (  posedge \AES.a1.S4_0.S_1.clk )
    begin
        case ( \AES.a1.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a1.S4_0.S_2.clk  = \AES.a1.S4_0.clk ;
    assign \AES.a1.S4_0.S_2.in  = \AES.a1.S4_0.in [15:8];
    assign \AES.a1.S4_0.k2  = \AES.a1.S4_0.S_2.out ;
    always @ (  posedge \AES.a1.S4_0.S_2.clk )
    begin
        case ( \AES.a1.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a1.S4_0.S_3.clk  = \AES.a1.S4_0.clk ;
    assign \AES.a1.S4_0.S_3.in  = \AES.a1.S4_0.in [7:0];
    assign \AES.a1.S4_0.k3  = \AES.a1.S4_0.S_3.out ;
    always @ (  posedge \AES.a1.S4_0.S_3.clk )
    begin
        case ( \AES.a1.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a1.S4_0.out  = { \AES.a1.S4_0.k0 , \AES.a1.S4_0.k1 , \AES.a1.S4_0.k2 , \AES.a1.S4_0.k3  };
    assign \AES.a1.k0b  = ( \AES.a1.k0a  ^ \AES.a1.k4a  );
    assign \AES.a1.k1b  = ( \AES.a1.k1a  ^ \AES.a1.k4a  );
    assign \AES.a1.k2b  = ( \AES.a1.k2a  ^ \AES.a1.k4a  );
    assign \AES.a1.k3b  = ( \AES.a1.k3a  ^ \AES.a1.k4a  );
    always @ (  posedge \AES.a1.clk )
    begin
    end
    assign \AES.a1.out_2  = { \AES.a1.k0b , \AES.a1.k1b , \AES.a1.k2b , \AES.a1.k3b  };
    assign \AES.a2.clk  = \AES.clk ;
    assign \AES.a2.in  = \AES.k1 ;
    assign \AES.a2.rcon  = \AES.k2 ;
    assign \AES.k1b  = \AES.a2.out_1 ;
    assign \AES.a2_rcon  = \AES.a2.out_2 ;
    assign \AES.a2.k0  = \AES.a2.in [127:96];
    assign \AES.a2.k1  = \AES.a2.in [95:64];
    assign \AES.a2.k2  = \AES.a2.in [63:32];
    assign \AES.a2.k3  = \AES.a2.in [31:0];
    assign \AES.a2.v0  = { ( \AES.a2.k0 [31:24] ^ \AES.a2.rcon  ), \AES.a2.k0 [23:0] };
    assign \AES.a2.v1  = ( \AES.a2.v0  ^ \AES.a2.k1  );
    assign \AES.a2.v2  = ( \AES.a2.v1  ^ \AES.a2.k2  );
    assign \AES.a2.v3  = ( \AES.a2.v2  ^ \AES.a2.k3  );
    always @ (  posedge \AES.a2.clk )
    begin
        \AES.a2.k0a  <= \AES.a2.v0 ;
        \AES.a2.k1a  <= \AES.a2.v1 ;
        \AES.a2.k2a  <= \AES.a2.v2 ;
        \AES.a2.k3a  <= \AES.a2.v3 ;
    end
    assign \AES.a2.S4_0.clk  = \AES.a2.clk ;
    assign \AES.a2.S4_0.in  = { \AES.a2.k3 [23:0], \AES.a2.k3 [31:24] };
    assign \AES.a2.k4a  = \AES.a2.S4_0.out ;
    assign \AES.a2.S4_0.S_0.clk  = \AES.a2.S4_0.clk ;
    assign \AES.a2.S4_0.S_0.in  = \AES.a2.S4_0.in [31:24];
    assign \AES.a2.S4_0.k0  = \AES.a2.S4_0.S_0.out ;
    always @ (  posedge \AES.a2.S4_0.S_0.clk )
    begin
        case ( \AES.a2.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a2.S4_0.S_1.clk  = \AES.a2.S4_0.clk ;
    assign \AES.a2.S4_0.S_1.in  = \AES.a2.S4_0.in [23:16];
    assign \AES.a2.S4_0.k1  = \AES.a2.S4_0.S_1.out ;
    always @ (  posedge \AES.a2.S4_0.S_1.clk )
    begin
        case ( \AES.a2.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a2.S4_0.S_2.clk  = \AES.a2.S4_0.clk ;
    assign \AES.a2.S4_0.S_2.in  = \AES.a2.S4_0.in [15:8];
    assign \AES.a2.S4_0.k2  = \AES.a2.S4_0.S_2.out ;
    always @ (  posedge \AES.a2.S4_0.S_2.clk )
    begin
        case ( \AES.a2.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a2.S4_0.S_3.clk  = \AES.a2.S4_0.clk ;
    assign \AES.a2.S4_0.S_3.in  = \AES.a2.S4_0.in [7:0];
    assign \AES.a2.S4_0.k3  = \AES.a2.S4_0.S_3.out ;
    always @ (  posedge \AES.a2.S4_0.S_3.clk )
    begin
        case ( \AES.a2.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a2.S4_0.out  = { \AES.a2.S4_0.k0 , \AES.a2.S4_0.k1 , \AES.a2.S4_0.k2 , \AES.a2.S4_0.k3  };
    assign \AES.a2.k0b  = ( \AES.a2.k0a  ^ \AES.a2.k4a  );
    assign \AES.a2.k1b  = ( \AES.a2.k1a  ^ \AES.a2.k4a  );
    assign \AES.a2.k2b  = ( \AES.a2.k2a  ^ \AES.a2.k4a  );
    assign \AES.a2.k3b  = ( \AES.a2.k3a  ^ \AES.a2.k4a  );
    always @ (  posedge \AES.a2.clk )
    begin
    end
    assign \AES.a2.out_2  = { \AES.a2.k0b , \AES.a2.k1b , \AES.a2.k2b , \AES.a2.k3b  };
    assign \AES.a3.clk  = \AES.clk ;
    assign \AES.a3.in  = \AES.k2 ;
    assign \AES.a3.rcon  = \AES.k3 ;
    assign \AES.k2b  = \AES.a3.out_1 ;
    assign \AES.a3_rcon  = \AES.a3.out_2 ;
    assign \AES.a3.k0  = \AES.a3.in [127:96];
    assign \AES.a3.k1  = \AES.a3.in [95:64];
    assign \AES.a3.k2  = \AES.a3.in [63:32];
    assign \AES.a3.k3  = \AES.a3.in [31:0];
    assign \AES.a3.v0  = { ( \AES.a3.k0 [31:24] ^ \AES.a3.rcon  ), \AES.a3.k0 [23:0] };
    assign \AES.a3.v1  = ( \AES.a3.v0  ^ \AES.a3.k1  );
    assign \AES.a3.v2  = ( \AES.a3.v1  ^ \AES.a3.k2  );
    assign \AES.a3.v3  = ( \AES.a3.v2  ^ \AES.a3.k3  );
    always @ (  posedge \AES.a3.clk )
    begin
        \AES.a3.k0a  <= \AES.a3.v0 ;
        \AES.a3.k1a  <= \AES.a3.v1 ;
        \AES.a3.k2a  <= \AES.a3.v2 ;
        \AES.a3.k3a  <= \AES.a3.v3 ;
    end
    assign \AES.a3.S4_0.clk  = \AES.a3.clk ;
    assign \AES.a3.S4_0.in  = { \AES.a3.k3 [23:0], \AES.a3.k3 [31:24] };
    assign \AES.a3.k4a  = \AES.a3.S4_0.out ;
    assign \AES.a3.S4_0.S_0.clk  = \AES.a3.S4_0.clk ;
    assign \AES.a3.S4_0.S_0.in  = \AES.a3.S4_0.in [31:24];
    assign \AES.a3.S4_0.k0  = \AES.a3.S4_0.S_0.out ;
    always @ (  posedge \AES.a3.S4_0.S_0.clk )
    begin
        case ( \AES.a3.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a3.S4_0.S_1.clk  = \AES.a3.S4_0.clk ;
    assign \AES.a3.S4_0.S_1.in  = \AES.a3.S4_0.in [23:16];
    assign \AES.a3.S4_0.k1  = \AES.a3.S4_0.S_1.out ;
    always @ (  posedge \AES.a3.S4_0.S_1.clk )
    begin
        case ( \AES.a3.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a3.S4_0.S_2.clk  = \AES.a3.S4_0.clk ;
    assign \AES.a3.S4_0.S_2.in  = \AES.a3.S4_0.in [15:8];
    assign \AES.a3.S4_0.k2  = \AES.a3.S4_0.S_2.out ;
    always @ (  posedge \AES.a3.S4_0.S_2.clk )
    begin
        case ( \AES.a3.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a3.S4_0.S_3.clk  = \AES.a3.S4_0.clk ;
    assign \AES.a3.S4_0.S_3.in  = \AES.a3.S4_0.in [7:0];
    assign \AES.a3.S4_0.k3  = \AES.a3.S4_0.S_3.out ;
    always @ (  posedge \AES.a3.S4_0.S_3.clk )
    begin
        case ( \AES.a3.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a3.S4_0.out  = { \AES.a3.S4_0.k0 , \AES.a3.S4_0.k1 , \AES.a3.S4_0.k2 , \AES.a3.S4_0.k3  };
    assign \AES.a3.k0b  = ( \AES.a3.k0a  ^ \AES.a3.k4a  );
    assign \AES.a3.k1b  = ( \AES.a3.k1a  ^ \AES.a3.k4a  );
    assign \AES.a3.k2b  = ( \AES.a3.k2a  ^ \AES.a3.k4a  );
    assign \AES.a3.k3b  = ( \AES.a3.k3a  ^ \AES.a3.k4a  );
    always @ (  posedge \AES.a3.clk )
    begin
    end
    assign \AES.a3.out_2  = { \AES.a3.k0b , \AES.a3.k1b , \AES.a3.k2b , \AES.a3.k3b  };
    assign \AES.a4.clk  = \AES.clk ;
    assign \AES.a4.in  = \AES.k3 ;
    assign \AES.a4.rcon  = \AES.k4 ;
    assign \AES.k3b  = \AES.a4.out_1 ;
    assign \AES.a4_rcon  = \AES.a4.out_2 ;
    assign \AES.a4.k0  = \AES.a4.in [127:96];
    assign \AES.a4.k1  = \AES.a4.in [95:64];
    assign \AES.a4.k2  = \AES.a4.in [63:32];
    assign \AES.a4.k3  = \AES.a4.in [31:0];
    assign \AES.a4.v0  = { ( \AES.a4.k0 [31:24] ^ \AES.a4.rcon  ), \AES.a4.k0 [23:0] };
    assign \AES.a4.v1  = ( \AES.a4.v0  ^ \AES.a4.k1  );
    assign \AES.a4.v2  = ( \AES.a4.v1  ^ \AES.a4.k2  );
    assign \AES.a4.v3  = ( \AES.a4.v2  ^ \AES.a4.k3  );
    always @ (  posedge \AES.a4.clk )
    begin
        \AES.a4.k0a  <= \AES.a4.v0 ;
        \AES.a4.k1a  <= \AES.a4.v1 ;
        \AES.a4.k2a  <= \AES.a4.v2 ;
        \AES.a4.k3a  <= \AES.a4.v3 ;
    end
    assign \AES.a4.S4_0.clk  = \AES.a4.clk ;
    assign \AES.a4.S4_0.in  = { \AES.a4.k3 [23:0], \AES.a4.k3 [31:24] };
    assign \AES.a4.k4a  = \AES.a4.S4_0.out ;
    assign \AES.a4.S4_0.S_0.clk  = \AES.a4.S4_0.clk ;
    assign \AES.a4.S4_0.S_0.in  = \AES.a4.S4_0.in [31:24];
    assign \AES.a4.S4_0.k0  = \AES.a4.S4_0.S_0.out ;
    always @ (  posedge \AES.a4.S4_0.S_0.clk )
    begin
        case ( \AES.a4.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a4.S4_0.S_1.clk  = \AES.a4.S4_0.clk ;
    assign \AES.a4.S4_0.S_1.in  = \AES.a4.S4_0.in [23:16];
    assign \AES.a4.S4_0.k1  = \AES.a4.S4_0.S_1.out ;
    always @ (  posedge \AES.a4.S4_0.S_1.clk )
    begin
        case ( \AES.a4.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a4.S4_0.S_2.clk  = \AES.a4.S4_0.clk ;
    assign \AES.a4.S4_0.S_2.in  = \AES.a4.S4_0.in [15:8];
    assign \AES.a4.S4_0.k2  = \AES.a4.S4_0.S_2.out ;
    always @ (  posedge \AES.a4.S4_0.S_2.clk )
    begin
        case ( \AES.a4.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a4.S4_0.S_3.clk  = \AES.a4.S4_0.clk ;
    assign \AES.a4.S4_0.S_3.in  = \AES.a4.S4_0.in [7:0];
    assign \AES.a4.S4_0.k3  = \AES.a4.S4_0.S_3.out ;
    always @ (  posedge \AES.a4.S4_0.S_3.clk )
    begin
        case ( \AES.a4.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a4.S4_0.out  = { \AES.a4.S4_0.k0 , \AES.a4.S4_0.k1 , \AES.a4.S4_0.k2 , \AES.a4.S4_0.k3  };
    assign \AES.a4.k0b  = ( \AES.a4.k0a  ^ \AES.a4.k4a  );
    assign \AES.a4.k1b  = ( \AES.a4.k1a  ^ \AES.a4.k4a  );
    assign \AES.a4.k2b  = ( \AES.a4.k2a  ^ \AES.a4.k4a  );
    assign \AES.a4.k3b  = ( \AES.a4.k3a  ^ \AES.a4.k4a  );
    always @ (  posedge \AES.a4.clk )
    begin
    end
    assign \AES.a4.out_2  = { \AES.a4.k0b , \AES.a4.k1b , \AES.a4.k2b , \AES.a4.k3b  };
    assign \AES.a5.clk  = \AES.clk ;
    assign \AES.a5.in  = \AES.k4 ;
    assign \AES.a5.rcon  = \AES.k5 ;
    assign \AES.k4b  = \AES.a5.out_1 ;
    assign \AES.a5_rcon  = \AES.a5.out_2 ;
    assign \AES.a5.k0  = \AES.a5.in [127:96];
    assign \AES.a5.k1  = \AES.a5.in [95:64];
    assign \AES.a5.k2  = \AES.a5.in [63:32];
    assign \AES.a5.k3  = \AES.a5.in [31:0];
    assign \AES.a5.v0  = { ( \AES.a5.k0 [31:24] ^ \AES.a5.rcon  ), \AES.a5.k0 [23:0] };
    assign \AES.a5.v1  = ( \AES.a5.v0  ^ \AES.a5.k1  );
    assign \AES.a5.v2  = ( \AES.a5.v1  ^ \AES.a5.k2  );
    assign \AES.a5.v3  = ( \AES.a5.v2  ^ \AES.a5.k3  );
    always @ (  posedge \AES.a5.clk )
    begin
        \AES.a5.k0a  <= \AES.a5.v0 ;
        \AES.a5.k1a  <= \AES.a5.v1 ;
        \AES.a5.k2a  <= \AES.a5.v2 ;
        \AES.a5.k3a  <= \AES.a5.v3 ;
    end
    assign \AES.a5.S4_0.clk  = \AES.a5.clk ;
    assign \AES.a5.S4_0.in  = { \AES.a5.k3 [23:0], \AES.a5.k3 [31:24] };
    assign \AES.a5.k4a  = \AES.a5.S4_0.out ;
    assign \AES.a5.S4_0.S_0.clk  = \AES.a5.S4_0.clk ;
    assign \AES.a5.S4_0.S_0.in  = \AES.a5.S4_0.in [31:24];
    assign \AES.a5.S4_0.k0  = \AES.a5.S4_0.S_0.out ;
    always @ (  posedge \AES.a5.S4_0.S_0.clk )
    begin
        case ( \AES.a5.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a5.S4_0.S_1.clk  = \AES.a5.S4_0.clk ;
    assign \AES.a5.S4_0.S_1.in  = \AES.a5.S4_0.in [23:16];
    assign \AES.a5.S4_0.k1  = \AES.a5.S4_0.S_1.out ;
    always @ (  posedge \AES.a5.S4_0.S_1.clk )
    begin
        case ( \AES.a5.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a5.S4_0.S_2.clk  = \AES.a5.S4_0.clk ;
    assign \AES.a5.S4_0.S_2.in  = \AES.a5.S4_0.in [15:8];
    assign \AES.a5.S4_0.k2  = \AES.a5.S4_0.S_2.out ;
    always @ (  posedge \AES.a5.S4_0.S_2.clk )
    begin
        case ( \AES.a5.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a5.S4_0.S_3.clk  = \AES.a5.S4_0.clk ;
    assign \AES.a5.S4_0.S_3.in  = \AES.a5.S4_0.in [7:0];
    assign \AES.a5.S4_0.k3  = \AES.a5.S4_0.S_3.out ;
    always @ (  posedge \AES.a5.S4_0.S_3.clk )
    begin
        case ( \AES.a5.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a5.S4_0.out  = { \AES.a5.S4_0.k0 , \AES.a5.S4_0.k1 , \AES.a5.S4_0.k2 , \AES.a5.S4_0.k3  };
    assign \AES.a5.k0b  = ( \AES.a5.k0a  ^ \AES.a5.k4a  );
    assign \AES.a5.k1b  = ( \AES.a5.k1a  ^ \AES.a5.k4a  );
    assign \AES.a5.k2b  = ( \AES.a5.k2a  ^ \AES.a5.k4a  );
    assign \AES.a5.k3b  = ( \AES.a5.k3a  ^ \AES.a5.k4a  );
    always @ (  posedge \AES.a5.clk )
    begin
    end
    assign \AES.a5.out_2  = { \AES.a5.k0b , \AES.a5.k1b , \AES.a5.k2b , \AES.a5.k3b  };
    assign \AES.a6.clk  = \AES.clk ;
    assign \AES.a6.in  = \AES.k5 ;
    assign \AES.a6.rcon  = \AES.k6 ;
    assign \AES.k5b  = \AES.a6.out_1 ;
    assign \AES.a6_rcon  = \AES.a6.out_2 ;
    assign \AES.a6.k0  = \AES.a6.in [127:96];
    assign \AES.a6.k1  = \AES.a6.in [95:64];
    assign \AES.a6.k2  = \AES.a6.in [63:32];
    assign \AES.a6.k3  = \AES.a6.in [31:0];
    assign \AES.a6.v0  = { ( \AES.a6.k0 [31:24] ^ \AES.a6.rcon  ), \AES.a6.k0 [23:0] };
    assign \AES.a6.v1  = ( \AES.a6.v0  ^ \AES.a6.k1  );
    assign \AES.a6.v2  = ( \AES.a6.v1  ^ \AES.a6.k2  );
    assign \AES.a6.v3  = ( \AES.a6.v2  ^ \AES.a6.k3  );
    always @ (  posedge \AES.a6.clk )
    begin
        \AES.a6.k0a  <= \AES.a6.v0 ;
        \AES.a6.k1a  <= \AES.a6.v1 ;
        \AES.a6.k2a  <= \AES.a6.v2 ;
        \AES.a6.k3a  <= \AES.a6.v3 ;
    end
    assign \AES.a6.S4_0.clk  = \AES.a6.clk ;
    assign \AES.a6.S4_0.in  = { \AES.a6.k3 [23:0], \AES.a6.k3 [31:24] };
    assign \AES.a6.k4a  = \AES.a6.S4_0.out ;
    assign \AES.a6.S4_0.S_0.clk  = \AES.a6.S4_0.clk ;
    assign \AES.a6.S4_0.S_0.in  = \AES.a6.S4_0.in [31:24];
    assign \AES.a6.S4_0.k0  = \AES.a6.S4_0.S_0.out ;
    always @ (  posedge \AES.a6.S4_0.S_0.clk )
    begin
        case ( \AES.a6.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a6.S4_0.S_1.clk  = \AES.a6.S4_0.clk ;
    assign \AES.a6.S4_0.S_1.in  = \AES.a6.S4_0.in [23:16];
    assign \AES.a6.S4_0.k1  = \AES.a6.S4_0.S_1.out ;
    always @ (  posedge \AES.a6.S4_0.S_1.clk )
    begin
        case ( \AES.a6.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a6.S4_0.S_2.clk  = \AES.a6.S4_0.clk ;
    assign \AES.a6.S4_0.S_2.in  = \AES.a6.S4_0.in [15:8];
    assign \AES.a6.S4_0.k2  = \AES.a6.S4_0.S_2.out ;
    always @ (  posedge \AES.a6.S4_0.S_2.clk )
    begin
        case ( \AES.a6.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a6.S4_0.S_3.clk  = \AES.a6.S4_0.clk ;
    assign \AES.a6.S4_0.S_3.in  = \AES.a6.S4_0.in [7:0];
    assign \AES.a6.S4_0.k3  = \AES.a6.S4_0.S_3.out ;
    always @ (  posedge \AES.a6.S4_0.S_3.clk )
    begin
        case ( \AES.a6.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a6.S4_0.out  = { \AES.a6.S4_0.k0 , \AES.a6.S4_0.k1 , \AES.a6.S4_0.k2 , \AES.a6.S4_0.k3  };
    assign \AES.a6.k0b  = ( \AES.a6.k0a  ^ \AES.a6.k4a  );
    assign \AES.a6.k1b  = ( \AES.a6.k1a  ^ \AES.a6.k4a  );
    assign \AES.a6.k2b  = ( \AES.a6.k2a  ^ \AES.a6.k4a  );
    assign \AES.a6.k3b  = ( \AES.a6.k3a  ^ \AES.a6.k4a  );
    always @ (  posedge \AES.a6.clk )
    begin
    end
    assign \AES.a6.out_2  = { \AES.a6.k0b , \AES.a6.k1b , \AES.a6.k2b , \AES.a6.k3b  };
    assign \AES.a7.clk  = \AES.clk ;
    assign \AES.a7.in  = \AES.k6 ;
    assign \AES.a7.rcon  = \AES.k7 ;
    assign \AES.k6b  = \AES.a7.out_1 ;
    assign \AES.a7_rcon  = \AES.a7.out_2 ;
    assign \AES.a7.k0  = \AES.a7.in [127:96];
    assign \AES.a7.k1  = \AES.a7.in [95:64];
    assign \AES.a7.k2  = \AES.a7.in [63:32];
    assign \AES.a7.k3  = \AES.a7.in [31:0];
    assign \AES.a7.v0  = { ( \AES.a7.k0 [31:24] ^ \AES.a7.rcon  ), \AES.a7.k0 [23:0] };
    assign \AES.a7.v1  = ( \AES.a7.v0  ^ \AES.a7.k1  );
    assign \AES.a7.v2  = ( \AES.a7.v1  ^ \AES.a7.k2  );
    assign \AES.a7.v3  = ( \AES.a7.v2  ^ \AES.a7.k3  );
    always @ (  posedge \AES.a7.clk )
    begin
        \AES.a7.k0a  <= \AES.a7.v0 ;
        \AES.a7.k1a  <= \AES.a7.v1 ;
        \AES.a7.k2a  <= \AES.a7.v2 ;
        \AES.a7.k3a  <= \AES.a7.v3 ;
    end
    assign \AES.a7.S4_0.clk  = \AES.a7.clk ;
    assign \AES.a7.S4_0.in  = { \AES.a7.k3 [23:0], \AES.a7.k3 [31:24] };
    assign \AES.a7.k4a  = \AES.a7.S4_0.out ;
    assign \AES.a7.S4_0.S_0.clk  = \AES.a7.S4_0.clk ;
    assign \AES.a7.S4_0.S_0.in  = \AES.a7.S4_0.in [31:24];
    assign \AES.a7.S4_0.k0  = \AES.a7.S4_0.S_0.out ;
    always @ (  posedge \AES.a7.S4_0.S_0.clk )
    begin
        case ( \AES.a7.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a7.S4_0.S_1.clk  = \AES.a7.S4_0.clk ;
    assign \AES.a7.S4_0.S_1.in  = \AES.a7.S4_0.in [23:16];
    assign \AES.a7.S4_0.k1  = \AES.a7.S4_0.S_1.out ;
    always @ (  posedge \AES.a7.S4_0.S_1.clk )
    begin
        case ( \AES.a7.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a7.S4_0.S_2.clk  = \AES.a7.S4_0.clk ;
    assign \AES.a7.S4_0.S_2.in  = \AES.a7.S4_0.in [15:8];
    assign \AES.a7.S4_0.k2  = \AES.a7.S4_0.S_2.out ;
    always @ (  posedge \AES.a7.S4_0.S_2.clk )
    begin
        case ( \AES.a7.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a7.S4_0.S_3.clk  = \AES.a7.S4_0.clk ;
    assign \AES.a7.S4_0.S_3.in  = \AES.a7.S4_0.in [7:0];
    assign \AES.a7.S4_0.k3  = \AES.a7.S4_0.S_3.out ;
    always @ (  posedge \AES.a7.S4_0.S_3.clk )
    begin
        case ( \AES.a7.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a7.S4_0.out  = { \AES.a7.S4_0.k0 , \AES.a7.S4_0.k1 , \AES.a7.S4_0.k2 , \AES.a7.S4_0.k3  };
    assign \AES.a7.k0b  = ( \AES.a7.k0a  ^ \AES.a7.k4a  );
    assign \AES.a7.k1b  = ( \AES.a7.k1a  ^ \AES.a7.k4a  );
    assign \AES.a7.k2b  = ( \AES.a7.k2a  ^ \AES.a7.k4a  );
    assign \AES.a7.k3b  = ( \AES.a7.k3a  ^ \AES.a7.k4a  );
    always @ (  posedge \AES.a7.clk )
    begin
    end
    assign \AES.a7.out_2  = { \AES.a7.k0b , \AES.a7.k1b , \AES.a7.k2b , \AES.a7.k3b  };
    assign \AES.a8.clk  = \AES.clk ;
    assign \AES.a8.in  = \AES.k7 ;
    assign \AES.a8.rcon  = \AES.k8 ;
    assign \AES.k7b  = \AES.a8.out_1 ;
    assign \AES.a8_rcon  = \AES.a8.out_2 ;
    assign \AES.a8.k0  = \AES.a8.in [127:96];
    assign \AES.a8.k1  = \AES.a8.in [95:64];
    assign \AES.a8.k2  = \AES.a8.in [63:32];
    assign \AES.a8.k3  = \AES.a8.in [31:0];
    assign \AES.a8.v0  = { ( \AES.a8.k0 [31:24] ^ \AES.a8.rcon  ), \AES.a8.k0 [23:0] };
    assign \AES.a8.v1  = ( \AES.a8.v0  ^ \AES.a8.k1  );
    assign \AES.a8.v2  = ( \AES.a8.v1  ^ \AES.a8.k2  );
    assign \AES.a8.v3  = ( \AES.a8.v2  ^ \AES.a8.k3  );
    always @ (  posedge \AES.a8.clk )
    begin
        \AES.a8.k0a  <= \AES.a8.v0 ;
        \AES.a8.k1a  <= \AES.a8.v1 ;
        \AES.a8.k2a  <= \AES.a8.v2 ;
        \AES.a8.k3a  <= \AES.a8.v3 ;
    end
    assign \AES.a8.S4_0.clk  = \AES.a8.clk ;
    assign \AES.a8.S4_0.in  = { \AES.a8.k3 [23:0], \AES.a8.k3 [31:24] };
    assign \AES.a8.k4a  = \AES.a8.S4_0.out ;
    assign \AES.a8.S4_0.S_0.clk  = \AES.a8.S4_0.clk ;
    assign \AES.a8.S4_0.S_0.in  = \AES.a8.S4_0.in [31:24];
    assign \AES.a8.S4_0.k0  = \AES.a8.S4_0.S_0.out ;
    always @ (  posedge \AES.a8.S4_0.S_0.clk )
    begin
        case ( \AES.a8.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a8.S4_0.S_1.clk  = \AES.a8.S4_0.clk ;
    assign \AES.a8.S4_0.S_1.in  = \AES.a8.S4_0.in [23:16];
    assign \AES.a8.S4_0.k1  = \AES.a8.S4_0.S_1.out ;
    always @ (  posedge \AES.a8.S4_0.S_1.clk )
    begin
        case ( \AES.a8.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a8.S4_0.S_2.clk  = \AES.a8.S4_0.clk ;
    assign \AES.a8.S4_0.S_2.in  = \AES.a8.S4_0.in [15:8];
    assign \AES.a8.S4_0.k2  = \AES.a8.S4_0.S_2.out ;
    always @ (  posedge \AES.a8.S4_0.S_2.clk )
    begin
        case ( \AES.a8.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a8.S4_0.S_3.clk  = \AES.a8.S4_0.clk ;
    assign \AES.a8.S4_0.S_3.in  = \AES.a8.S4_0.in [7:0];
    assign \AES.a8.S4_0.k3  = \AES.a8.S4_0.S_3.out ;
    always @ (  posedge \AES.a8.S4_0.S_3.clk )
    begin
        case ( \AES.a8.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a8.S4_0.out  = { \AES.a8.S4_0.k0 , \AES.a8.S4_0.k1 , \AES.a8.S4_0.k2 , \AES.a8.S4_0.k3  };
    assign \AES.a8.k0b  = ( \AES.a8.k0a  ^ \AES.a8.k4a  );
    assign \AES.a8.k1b  = ( \AES.a8.k1a  ^ \AES.a8.k4a  );
    assign \AES.a8.k2b  = ( \AES.a8.k2a  ^ \AES.a8.k4a  );
    assign \AES.a8.k3b  = ( \AES.a8.k3a  ^ \AES.a8.k4a  );
    always @ (  posedge \AES.a8.clk )
    begin
    end
    assign \AES.a8.out_2  = { \AES.a8.k0b , \AES.a8.k1b , \AES.a8.k2b , \AES.a8.k3b  };
    assign \AES.a9.clk  = \AES.clk ;
    assign \AES.a9.in  = \AES.k8 ;
    assign \AES.a9.rcon  = \AES.k9 ;
    assign \AES.k8b  = \AES.a9.out_1 ;
    assign \AES.a9_rcon  = \AES.a9.out_2 ;
    assign \AES.a9.k0  = \AES.a9.in [127:96];
    assign \AES.a9.k1  = \AES.a9.in [95:64];
    assign \AES.a9.k2  = \AES.a9.in [63:32];
    assign \AES.a9.k3  = \AES.a9.in [31:0];
    assign \AES.a9.v0  = { ( \AES.a9.k0 [31:24] ^ \AES.a9.rcon  ), \AES.a9.k0 [23:0] };
    assign \AES.a9.v1  = ( \AES.a9.v0  ^ \AES.a9.k1  );
    assign \AES.a9.v2  = ( \AES.a9.v1  ^ \AES.a9.k2  );
    assign \AES.a9.v3  = ( \AES.a9.v2  ^ \AES.a9.k3  );
    always @ (  posedge \AES.a9.clk )
    begin
        \AES.a9.k0a  <= \AES.a9.v0 ;
        \AES.a9.k1a  <= \AES.a9.v1 ;
        \AES.a9.k2a  <= \AES.a9.v2 ;
        \AES.a9.k3a  <= \AES.a9.v3 ;
    end
    assign \AES.a9.S4_0.clk  = \AES.a9.clk ;
    assign \AES.a9.S4_0.in  = { \AES.a9.k3 [23:0], \AES.a9.k3 [31:24] };
    assign \AES.a9.k4a  = \AES.a9.S4_0.out ;
    assign \AES.a9.S4_0.S_0.clk  = \AES.a9.S4_0.clk ;
    assign \AES.a9.S4_0.S_0.in  = \AES.a9.S4_0.in [31:24];
    assign \AES.a9.S4_0.k0  = \AES.a9.S4_0.S_0.out ;
    always @ (  posedge \AES.a9.S4_0.S_0.clk )
    begin
        case ( \AES.a9.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a9.S4_0.S_1.clk  = \AES.a9.S4_0.clk ;
    assign \AES.a9.S4_0.S_1.in  = \AES.a9.S4_0.in [23:16];
    assign \AES.a9.S4_0.k1  = \AES.a9.S4_0.S_1.out ;
    always @ (  posedge \AES.a9.S4_0.S_1.clk )
    begin
        case ( \AES.a9.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a9.S4_0.S_2.clk  = \AES.a9.S4_0.clk ;
    assign \AES.a9.S4_0.S_2.in  = \AES.a9.S4_0.in [15:8];
    assign \AES.a9.S4_0.k2  = \AES.a9.S4_0.S_2.out ;
    always @ (  posedge \AES.a9.S4_0.S_2.clk )
    begin
        case ( \AES.a9.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a9.S4_0.S_3.clk  = \AES.a9.S4_0.clk ;
    assign \AES.a9.S4_0.S_3.in  = \AES.a9.S4_0.in [7:0];
    assign \AES.a9.S4_0.k3  = \AES.a9.S4_0.S_3.out ;
    always @ (  posedge \AES.a9.S4_0.S_3.clk )
    begin
        case ( \AES.a9.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a9.S4_0.out  = { \AES.a9.S4_0.k0 , \AES.a9.S4_0.k1 , \AES.a9.S4_0.k2 , \AES.a9.S4_0.k3  };
    assign \AES.a9.k0b  = ( \AES.a9.k0a  ^ \AES.a9.k4a  );
    assign \AES.a9.k1b  = ( \AES.a9.k1a  ^ \AES.a9.k4a  );
    assign \AES.a9.k2b  = ( \AES.a9.k2a  ^ \AES.a9.k4a  );
    assign \AES.a9.k3b  = ( \AES.a9.k3a  ^ \AES.a9.k4a  );
    always @ (  posedge \AES.a9.clk )
    begin
    end
    assign \AES.a9.out_2  = { \AES.a9.k0b , \AES.a9.k1b , \AES.a9.k2b , \AES.a9.k3b  };
    assign \AES.a10.clk  = \AES.clk ;
    assign \AES.a10.in  = \AES.k9 ;
    assign \AES.a10.rcon  = \AES.k10 ;
    assign \AES.k9b  = \AES.a10.out_1 ;
    assign \AES.a10_rcon  = \AES.a10.out_2 ;
    assign \AES.a10.k0  = \AES.a10.in [127:96];
    assign \AES.a10.k1  = \AES.a10.in [95:64];
    assign \AES.a10.k2  = \AES.a10.in [63:32];
    assign \AES.a10.k3  = \AES.a10.in [31:0];
    assign \AES.a10.v0  = { ( \AES.a10.k0 [31:24] ^ \AES.a10.rcon  ), \AES.a10.k0 [23:0] };
    assign \AES.a10.v1  = ( \AES.a10.v0  ^ \AES.a10.k1  );
    assign \AES.a10.v2  = ( \AES.a10.v1  ^ \AES.a10.k2  );
    assign \AES.a10.v3  = ( \AES.a10.v2  ^ \AES.a10.k3  );
    always @ (  posedge \AES.a10.clk )
    begin
        \AES.a10.k0a  <= \AES.a10.v0 ;
        \AES.a10.k1a  <= \AES.a10.v1 ;
        \AES.a10.k2a  <= \AES.a10.v2 ;
        \AES.a10.k3a  <= \AES.a10.v3 ;
    end
    assign \AES.a10.S4_0.clk  = \AES.a10.clk ;
    assign \AES.a10.S4_0.in  = { \AES.a10.k3 [23:0], \AES.a10.k3 [31:24] };
    assign \AES.a10.k4a  = \AES.a10.S4_0.out ;
    assign \AES.a10.S4_0.S_0.clk  = \AES.a10.S4_0.clk ;
    assign \AES.a10.S4_0.S_0.in  = \AES.a10.S4_0.in [31:24];
    assign \AES.a10.S4_0.k0  = \AES.a10.S4_0.S_0.out ;
    always @ (  posedge \AES.a10.S4_0.S_0.clk )
    begin
        case ( \AES.a10.S4_0.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a10.S4_0.S_1.clk  = \AES.a10.S4_0.clk ;
    assign \AES.a10.S4_0.S_1.in  = \AES.a10.S4_0.in [23:16];
    assign \AES.a10.S4_0.k1  = \AES.a10.S4_0.S_1.out ;
    always @ (  posedge \AES.a10.S4_0.S_1.clk )
    begin
        case ( \AES.a10.S4_0.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a10.S4_0.S_2.clk  = \AES.a10.S4_0.clk ;
    assign \AES.a10.S4_0.S_2.in  = \AES.a10.S4_0.in [15:8];
    assign \AES.a10.S4_0.k2  = \AES.a10.S4_0.S_2.out ;
    always @ (  posedge \AES.a10.S4_0.S_2.clk )
    begin
        case ( \AES.a10.S4_0.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a10.S4_0.S_3.clk  = \AES.a10.S4_0.clk ;
    assign \AES.a10.S4_0.S_3.in  = \AES.a10.S4_0.in [7:0];
    assign \AES.a10.S4_0.k3  = \AES.a10.S4_0.S_3.out ;
    always @ (  posedge \AES.a10.S4_0.S_3.clk )
    begin
        case ( \AES.a10.S4_0.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.a10.S4_0.out  = { \AES.a10.S4_0.k0 , \AES.a10.S4_0.k1 , \AES.a10.S4_0.k2 , \AES.a10.S4_0.k3  };
    assign \AES.a10.k0b  = ( \AES.a10.k0a  ^ \AES.a10.k4a  );
    assign \AES.a10.k1b  = ( \AES.a10.k1a  ^ \AES.a10.k4a  );
    assign \AES.a10.k2b  = ( \AES.a10.k2a  ^ \AES.a10.k4a  );
    assign \AES.a10.k3b  = ( \AES.a10.k3a  ^ \AES.a10.k4a  );
    always @ (  posedge \AES.a10.clk )
    begin
    end
    assign \AES.a10.out_2  = { \AES.a10.k0b , \AES.a10.k1b , \AES.a10.k2b , \AES.a10.k3b  };
    assign \AES.r1.clk  = \AES.clk ;
    assign \AES.r1.state_in  = \AES.s0 ;
    assign \AES.r1.key  = \AES.k0b ;
    assign \AES.s1  = \AES.r1.state_out ;
    assign \AES.r1.k0  = \AES.r1.key [127:96];
    assign \AES.r1.k1  = \AES.r1.key [95:64];
    assign \AES.r1.k2  = \AES.r1.key [63:32];
    assign \AES.r1.k3  = \AES.r1.key [31:0];
    assign \AES.r1.s0  = \AES.r1.state_in [127:96];
    assign \AES.r1.s1  = \AES.r1.state_in [95:64];
    assign \AES.r1.s2  = \AES.r1.state_in [63:32];
    assign \AES.r1.s3  = \AES.r1.state_in [31:0];
    assign \AES.r1.t0.clk  = \AES.r1.clk ;
    assign \AES.r1.t0.state  = \AES.r1.s0 ;
    assign \AES.r1.p00  = \AES.r1.t0.p0 ;
    assign \AES.r1.p01  = \AES.r1.t0.p1 ;
    assign \AES.r1.p02  = \AES.r1.t0.p2 ;
    assign \AES.r1.p03  = \AES.r1.t0.p3 ;
    assign \AES.r1.t0.p0  = { \AES.r1.t0.k0 [7:0], \AES.r1.t0.k0 [31:8] };
    assign \AES.r1.t0.p1  = { \AES.r1.t0.k1 [15:0], \AES.r1.t0.k1 [31:16] };
    assign \AES.r1.t0.p2  = { \AES.r1.t0.k2 [23:0], \AES.r1.t0.k2 [31:24] };
    assign \AES.r1.t0.b0  = \AES.r1.t0.state [31:24];
    assign \AES.r1.t0.b1  = \AES.r1.t0.state [23:16];
    assign \AES.r1.t0.b2  = \AES.r1.t0.state [15:8];
    assign \AES.r1.t0.b3  = \AES.r1.t0.state [7:0];
    assign \AES.r1.t0.t0.clk  = \AES.r1.t0.clk ;
    assign \AES.r1.t0.t0.in  = \AES.r1.t0.b0 ;
    assign \AES.r1.t0.k0  = \AES.r1.t0.t0.out ;
    assign \AES.r1.t0.t0.s0.clk  = \AES.r1.t0.t0.clk ;
    assign \AES.r1.t0.t0.s0.in  = \AES.r1.t0.t0.in ;
    assign \AES.r1.t0.t0.k0  = \AES.r1.t0.t0.s0.out ;
    always @ (  posedge \AES.r1.t0.t0.s0.clk )
    begin
        case ( \AES.r1.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t0.s4.clk  = \AES.r1.t0.t0.clk ;
    assign \AES.r1.t0.t0.s4.in  = \AES.r1.t0.t0.in ;
    assign \AES.r1.t0.t0.k1  = \AES.r1.t0.t0.s4.out ;
    always @ (  posedge \AES.r1.t0.t0.s4.clk )
    begin
        case ( \AES.r1.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t0.out  = { \AES.r1.t0.t0.k0 , \AES.r1.t0.t0.k0 , ( \AES.r1.t0.t0.k0  ^ \AES.r1.t0.t0.k1  ), \AES.r1.t0.t0.k1  };
    assign \AES.r1.t0.t1.clk  = \AES.r1.t0.clk ;
    assign \AES.r1.t0.t1.in  = \AES.r1.t0.b1 ;
    assign \AES.r1.t0.k1  = \AES.r1.t0.t1.out ;
    assign \AES.r1.t0.t1.s0.clk  = \AES.r1.t0.t1.clk ;
    assign \AES.r1.t0.t1.s0.in  = \AES.r1.t0.t1.in ;
    assign \AES.r1.t0.t1.k0  = \AES.r1.t0.t1.s0.out ;
    always @ (  posedge \AES.r1.t0.t1.s0.clk )
    begin
        case ( \AES.r1.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t1.s4.clk  = \AES.r1.t0.t1.clk ;
    assign \AES.r1.t0.t1.s4.in  = \AES.r1.t0.t1.in ;
    assign \AES.r1.t0.t1.k1  = \AES.r1.t0.t1.s4.out ;
    always @ (  posedge \AES.r1.t0.t1.s4.clk )
    begin
        case ( \AES.r1.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t1.out  = { \AES.r1.t0.t1.k0 , \AES.r1.t0.t1.k0 , ( \AES.r1.t0.t1.k0  ^ \AES.r1.t0.t1.k1  ), \AES.r1.t0.t1.k1  };
    assign \AES.r1.t0.t2.clk  = \AES.r1.t0.clk ;
    assign \AES.r1.t0.t2.in  = \AES.r1.t0.b2 ;
    assign \AES.r1.t0.k2  = \AES.r1.t0.t2.out ;
    assign \AES.r1.t0.t2.s0.clk  = \AES.r1.t0.t2.clk ;
    assign \AES.r1.t0.t2.s0.in  = \AES.r1.t0.t2.in ;
    assign \AES.r1.t0.t2.k0  = \AES.r1.t0.t2.s0.out ;
    always @ (  posedge \AES.r1.t0.t2.s0.clk )
    begin
        case ( \AES.r1.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t2.s4.clk  = \AES.r1.t0.t2.clk ;
    assign \AES.r1.t0.t2.s4.in  = \AES.r1.t0.t2.in ;
    assign \AES.r1.t0.t2.k1  = \AES.r1.t0.t2.s4.out ;
    always @ (  posedge \AES.r1.t0.t2.s4.clk )
    begin
        case ( \AES.r1.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t2.out  = { \AES.r1.t0.t2.k0 , \AES.r1.t0.t2.k0 , ( \AES.r1.t0.t2.k0  ^ \AES.r1.t0.t2.k1  ), \AES.r1.t0.t2.k1  };
    assign \AES.r1.t0.t3.clk  = \AES.r1.t0.clk ;
    assign \AES.r1.t0.t3.in  = \AES.r1.t0.b3 ;
    assign \AES.r1.t0.p3  = \AES.r1.t0.t3.out ;
    assign \AES.r1.t0.t3.s0.clk  = \AES.r1.t0.t3.clk ;
    assign \AES.r1.t0.t3.s0.in  = \AES.r1.t0.t3.in ;
    assign \AES.r1.t0.t3.k0  = \AES.r1.t0.t3.s0.out ;
    always @ (  posedge \AES.r1.t0.t3.s0.clk )
    begin
        case ( \AES.r1.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t3.s4.clk  = \AES.r1.t0.t3.clk ;
    assign \AES.r1.t0.t3.s4.in  = \AES.r1.t0.t3.in ;
    assign \AES.r1.t0.t3.k1  = \AES.r1.t0.t3.s4.out ;
    always @ (  posedge \AES.r1.t0.t3.s4.clk )
    begin
        case ( \AES.r1.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t0.t3.out  = { \AES.r1.t0.t3.k0 , \AES.r1.t0.t3.k0 , ( \AES.r1.t0.t3.k0  ^ \AES.r1.t0.t3.k1  ), \AES.r1.t0.t3.k1  };
    assign \AES.r1.t1.clk  = \AES.r1.clk ;
    assign \AES.r1.t1.state  = \AES.r1.s1 ;
    assign \AES.r1.p10  = \AES.r1.t1.p0 ;
    assign \AES.r1.p11  = \AES.r1.t1.p1 ;
    assign \AES.r1.p12  = \AES.r1.t1.p2 ;
    assign \AES.r1.p13  = \AES.r1.t1.p3 ;
    assign \AES.r1.t1.p0  = { \AES.r1.t1.k0 [7:0], \AES.r1.t1.k0 [31:8] };
    assign \AES.r1.t1.p1  = { \AES.r1.t1.k1 [15:0], \AES.r1.t1.k1 [31:16] };
    assign \AES.r1.t1.p2  = { \AES.r1.t1.k2 [23:0], \AES.r1.t1.k2 [31:24] };
    assign \AES.r1.t1.b0  = \AES.r1.t1.state [31:24];
    assign \AES.r1.t1.b1  = \AES.r1.t1.state [23:16];
    assign \AES.r1.t1.b2  = \AES.r1.t1.state [15:8];
    assign \AES.r1.t1.b3  = \AES.r1.t1.state [7:0];
    assign \AES.r1.t1.t0.clk  = \AES.r1.t1.clk ;
    assign \AES.r1.t1.t0.in  = \AES.r1.t1.b0 ;
    assign \AES.r1.t1.k0  = \AES.r1.t1.t0.out ;
    assign \AES.r1.t1.t0.s0.clk  = \AES.r1.t1.t0.clk ;
    assign \AES.r1.t1.t0.s0.in  = \AES.r1.t1.t0.in ;
    assign \AES.r1.t1.t0.k0  = \AES.r1.t1.t0.s0.out ;
    always @ (  posedge \AES.r1.t1.t0.s0.clk )
    begin
        case ( \AES.r1.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t0.s4.clk  = \AES.r1.t1.t0.clk ;
    assign \AES.r1.t1.t0.s4.in  = \AES.r1.t1.t0.in ;
    assign \AES.r1.t1.t0.k1  = \AES.r1.t1.t0.s4.out ;
    always @ (  posedge \AES.r1.t1.t0.s4.clk )
    begin
        case ( \AES.r1.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t0.out  = { \AES.r1.t1.t0.k0 , \AES.r1.t1.t0.k0 , ( \AES.r1.t1.t0.k0  ^ \AES.r1.t1.t0.k1  ), \AES.r1.t1.t0.k1  };
    assign \AES.r1.t1.t1.clk  = \AES.r1.t1.clk ;
    assign \AES.r1.t1.t1.in  = \AES.r1.t1.b1 ;
    assign \AES.r1.t1.k1  = \AES.r1.t1.t1.out ;
    assign \AES.r1.t1.t1.s0.clk  = \AES.r1.t1.t1.clk ;
    assign \AES.r1.t1.t1.s0.in  = \AES.r1.t1.t1.in ;
    assign \AES.r1.t1.t1.k0  = \AES.r1.t1.t1.s0.out ;
    always @ (  posedge \AES.r1.t1.t1.s0.clk )
    begin
        case ( \AES.r1.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t1.s4.clk  = \AES.r1.t1.t1.clk ;
    assign \AES.r1.t1.t1.s4.in  = \AES.r1.t1.t1.in ;
    assign \AES.r1.t1.t1.k1  = \AES.r1.t1.t1.s4.out ;
    always @ (  posedge \AES.r1.t1.t1.s4.clk )
    begin
        case ( \AES.r1.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t1.out  = { \AES.r1.t1.t1.k0 , \AES.r1.t1.t1.k0 , ( \AES.r1.t1.t1.k0  ^ \AES.r1.t1.t1.k1  ), \AES.r1.t1.t1.k1  };
    assign \AES.r1.t1.t2.clk  = \AES.r1.t1.clk ;
    assign \AES.r1.t1.t2.in  = \AES.r1.t1.b2 ;
    assign \AES.r1.t1.k2  = \AES.r1.t1.t2.out ;
    assign \AES.r1.t1.t2.s0.clk  = \AES.r1.t1.t2.clk ;
    assign \AES.r1.t1.t2.s0.in  = \AES.r1.t1.t2.in ;
    assign \AES.r1.t1.t2.k0  = \AES.r1.t1.t2.s0.out ;
    always @ (  posedge \AES.r1.t1.t2.s0.clk )
    begin
        case ( \AES.r1.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t2.s4.clk  = \AES.r1.t1.t2.clk ;
    assign \AES.r1.t1.t2.s4.in  = \AES.r1.t1.t2.in ;
    assign \AES.r1.t1.t2.k1  = \AES.r1.t1.t2.s4.out ;
    always @ (  posedge \AES.r1.t1.t2.s4.clk )
    begin
        case ( \AES.r1.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t2.out  = { \AES.r1.t1.t2.k0 , \AES.r1.t1.t2.k0 , ( \AES.r1.t1.t2.k0  ^ \AES.r1.t1.t2.k1  ), \AES.r1.t1.t2.k1  };
    assign \AES.r1.t1.t3.clk  = \AES.r1.t1.clk ;
    assign \AES.r1.t1.t3.in  = \AES.r1.t1.b3 ;
    assign \AES.r1.t1.p3  = \AES.r1.t1.t3.out ;
    assign \AES.r1.t1.t3.s0.clk  = \AES.r1.t1.t3.clk ;
    assign \AES.r1.t1.t3.s0.in  = \AES.r1.t1.t3.in ;
    assign \AES.r1.t1.t3.k0  = \AES.r1.t1.t3.s0.out ;
    always @ (  posedge \AES.r1.t1.t3.s0.clk )
    begin
        case ( \AES.r1.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t3.s4.clk  = \AES.r1.t1.t3.clk ;
    assign \AES.r1.t1.t3.s4.in  = \AES.r1.t1.t3.in ;
    assign \AES.r1.t1.t3.k1  = \AES.r1.t1.t3.s4.out ;
    always @ (  posedge \AES.r1.t1.t3.s4.clk )
    begin
        case ( \AES.r1.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t1.t3.out  = { \AES.r1.t1.t3.k0 , \AES.r1.t1.t3.k0 , ( \AES.r1.t1.t3.k0  ^ \AES.r1.t1.t3.k1  ), \AES.r1.t1.t3.k1  };
    assign \AES.r1.t2.clk  = \AES.r1.clk ;
    assign \AES.r1.t2.state  = \AES.r1.s2 ;
    assign \AES.r1.p20  = \AES.r1.t2.p0 ;
    assign \AES.r1.p21  = \AES.r1.t2.p1 ;
    assign \AES.r1.p22  = \AES.r1.t2.p2 ;
    assign \AES.r1.p23  = \AES.r1.t2.p3 ;
    assign \AES.r1.t2.p0  = { \AES.r1.t2.k0 [7:0], \AES.r1.t2.k0 [31:8] };
    assign \AES.r1.t2.p1  = { \AES.r1.t2.k1 [15:0], \AES.r1.t2.k1 [31:16] };
    assign \AES.r1.t2.p2  = { \AES.r1.t2.k2 [23:0], \AES.r1.t2.k2 [31:24] };
    assign \AES.r1.t2.b0  = \AES.r1.t2.state [31:24];
    assign \AES.r1.t2.b1  = \AES.r1.t2.state [23:16];
    assign \AES.r1.t2.b2  = \AES.r1.t2.state [15:8];
    assign \AES.r1.t2.b3  = \AES.r1.t2.state [7:0];
    assign \AES.r1.t2.t0.clk  = \AES.r1.t2.clk ;
    assign \AES.r1.t2.t0.in  = \AES.r1.t2.b0 ;
    assign \AES.r1.t2.k0  = \AES.r1.t2.t0.out ;
    assign \AES.r1.t2.t0.s0.clk  = \AES.r1.t2.t0.clk ;
    assign \AES.r1.t2.t0.s0.in  = \AES.r1.t2.t0.in ;
    assign \AES.r1.t2.t0.k0  = \AES.r1.t2.t0.s0.out ;
    always @ (  posedge \AES.r1.t2.t0.s0.clk )
    begin
        case ( \AES.r1.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t0.s4.clk  = \AES.r1.t2.t0.clk ;
    assign \AES.r1.t2.t0.s4.in  = \AES.r1.t2.t0.in ;
    assign \AES.r1.t2.t0.k1  = \AES.r1.t2.t0.s4.out ;
    always @ (  posedge \AES.r1.t2.t0.s4.clk )
    begin
        case ( \AES.r1.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t0.out  = { \AES.r1.t2.t0.k0 , \AES.r1.t2.t0.k0 , ( \AES.r1.t2.t0.k0  ^ \AES.r1.t2.t0.k1  ), \AES.r1.t2.t0.k1  };
    assign \AES.r1.t2.t1.clk  = \AES.r1.t2.clk ;
    assign \AES.r1.t2.t1.in  = \AES.r1.t2.b1 ;
    assign \AES.r1.t2.k1  = \AES.r1.t2.t1.out ;
    assign \AES.r1.t2.t1.s0.clk  = \AES.r1.t2.t1.clk ;
    assign \AES.r1.t2.t1.s0.in  = \AES.r1.t2.t1.in ;
    assign \AES.r1.t2.t1.k0  = \AES.r1.t2.t1.s0.out ;
    always @ (  posedge \AES.r1.t2.t1.s0.clk )
    begin
        case ( \AES.r1.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t1.s4.clk  = \AES.r1.t2.t1.clk ;
    assign \AES.r1.t2.t1.s4.in  = \AES.r1.t2.t1.in ;
    assign \AES.r1.t2.t1.k1  = \AES.r1.t2.t1.s4.out ;
    always @ (  posedge \AES.r1.t2.t1.s4.clk )
    begin
        case ( \AES.r1.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t1.out  = { \AES.r1.t2.t1.k0 , \AES.r1.t2.t1.k0 , ( \AES.r1.t2.t1.k0  ^ \AES.r1.t2.t1.k1  ), \AES.r1.t2.t1.k1  };
    assign \AES.r1.t2.t2.clk  = \AES.r1.t2.clk ;
    assign \AES.r1.t2.t2.in  = \AES.r1.t2.b2 ;
    assign \AES.r1.t2.k2  = \AES.r1.t2.t2.out ;
    assign \AES.r1.t2.t2.s0.clk  = \AES.r1.t2.t2.clk ;
    assign \AES.r1.t2.t2.s0.in  = \AES.r1.t2.t2.in ;
    assign \AES.r1.t2.t2.k0  = \AES.r1.t2.t2.s0.out ;
    always @ (  posedge \AES.r1.t2.t2.s0.clk )
    begin
        case ( \AES.r1.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t2.s4.clk  = \AES.r1.t2.t2.clk ;
    assign \AES.r1.t2.t2.s4.in  = \AES.r1.t2.t2.in ;
    assign \AES.r1.t2.t2.k1  = \AES.r1.t2.t2.s4.out ;
    always @ (  posedge \AES.r1.t2.t2.s4.clk )
    begin
        case ( \AES.r1.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t2.out  = { \AES.r1.t2.t2.k0 , \AES.r1.t2.t2.k0 , ( \AES.r1.t2.t2.k0  ^ \AES.r1.t2.t2.k1  ), \AES.r1.t2.t2.k1  };
    assign \AES.r1.t2.t3.clk  = \AES.r1.t2.clk ;
    assign \AES.r1.t2.t3.in  = \AES.r1.t2.b3 ;
    assign \AES.r1.t2.p3  = \AES.r1.t2.t3.out ;
    assign \AES.r1.t2.t3.s0.clk  = \AES.r1.t2.t3.clk ;
    assign \AES.r1.t2.t3.s0.in  = \AES.r1.t2.t3.in ;
    assign \AES.r1.t2.t3.k0  = \AES.r1.t2.t3.s0.out ;
    always @ (  posedge \AES.r1.t2.t3.s0.clk )
    begin
        case ( \AES.r1.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t3.s4.clk  = \AES.r1.t2.t3.clk ;
    assign \AES.r1.t2.t3.s4.in  = \AES.r1.t2.t3.in ;
    assign \AES.r1.t2.t3.k1  = \AES.r1.t2.t3.s4.out ;
    always @ (  posedge \AES.r1.t2.t3.s4.clk )
    begin
        case ( \AES.r1.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t2.t3.out  = { \AES.r1.t2.t3.k0 , \AES.r1.t2.t3.k0 , ( \AES.r1.t2.t3.k0  ^ \AES.r1.t2.t3.k1  ), \AES.r1.t2.t3.k1  };
    assign \AES.r1.t3.clk  = \AES.r1.clk ;
    assign \AES.r1.t3.state  = \AES.r1.s3 ;
    assign \AES.r1.p30  = \AES.r1.t3.p0 ;
    assign \AES.r1.p31  = \AES.r1.t3.p1 ;
    assign \AES.r1.p32  = \AES.r1.t3.p2 ;
    assign \AES.r1.p33  = \AES.r1.t3.p3 ;
    assign \AES.r1.t3.p0  = { \AES.r1.t3.k0 [7:0], \AES.r1.t3.k0 [31:8] };
    assign \AES.r1.t3.p1  = { \AES.r1.t3.k1 [15:0], \AES.r1.t3.k1 [31:16] };
    assign \AES.r1.t3.p2  = { \AES.r1.t3.k2 [23:0], \AES.r1.t3.k2 [31:24] };
    assign \AES.r1.t3.b0  = \AES.r1.t3.state [31:24];
    assign \AES.r1.t3.b1  = \AES.r1.t3.state [23:16];
    assign \AES.r1.t3.b2  = \AES.r1.t3.state [15:8];
    assign \AES.r1.t3.b3  = \AES.r1.t3.state [7:0];
    assign \AES.r1.t3.t0.clk  = \AES.r1.t3.clk ;
    assign \AES.r1.t3.t0.in  = \AES.r1.t3.b0 ;
    assign \AES.r1.t3.k0  = \AES.r1.t3.t0.out ;
    assign \AES.r1.t3.t0.s0.clk  = \AES.r1.t3.t0.clk ;
    assign \AES.r1.t3.t0.s0.in  = \AES.r1.t3.t0.in ;
    assign \AES.r1.t3.t0.k0  = \AES.r1.t3.t0.s0.out ;
    always @ (  posedge \AES.r1.t3.t0.s0.clk )
    begin
        case ( \AES.r1.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t0.s4.clk  = \AES.r1.t3.t0.clk ;
    assign \AES.r1.t3.t0.s4.in  = \AES.r1.t3.t0.in ;
    assign \AES.r1.t3.t0.k1  = \AES.r1.t3.t0.s4.out ;
    always @ (  posedge \AES.r1.t3.t0.s4.clk )
    begin
        case ( \AES.r1.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t0.out  = { \AES.r1.t3.t0.k0 , \AES.r1.t3.t0.k0 , ( \AES.r1.t3.t0.k0  ^ \AES.r1.t3.t0.k1  ), \AES.r1.t3.t0.k1  };
    assign \AES.r1.t3.t1.clk  = \AES.r1.t3.clk ;
    assign \AES.r1.t3.t1.in  = \AES.r1.t3.b1 ;
    assign \AES.r1.t3.k1  = \AES.r1.t3.t1.out ;
    assign \AES.r1.t3.t1.s0.clk  = \AES.r1.t3.t1.clk ;
    assign \AES.r1.t3.t1.s0.in  = \AES.r1.t3.t1.in ;
    assign \AES.r1.t3.t1.k0  = \AES.r1.t3.t1.s0.out ;
    always @ (  posedge \AES.r1.t3.t1.s0.clk )
    begin
        case ( \AES.r1.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t1.s4.clk  = \AES.r1.t3.t1.clk ;
    assign \AES.r1.t3.t1.s4.in  = \AES.r1.t3.t1.in ;
    assign \AES.r1.t3.t1.k1  = \AES.r1.t3.t1.s4.out ;
    always @ (  posedge \AES.r1.t3.t1.s4.clk )
    begin
        case ( \AES.r1.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t1.out  = { \AES.r1.t3.t1.k0 , \AES.r1.t3.t1.k0 , ( \AES.r1.t3.t1.k0  ^ \AES.r1.t3.t1.k1  ), \AES.r1.t3.t1.k1  };
    assign \AES.r1.t3.t2.clk  = \AES.r1.t3.clk ;
    assign \AES.r1.t3.t2.in  = \AES.r1.t3.b2 ;
    assign \AES.r1.t3.k2  = \AES.r1.t3.t2.out ;
    assign \AES.r1.t3.t2.s0.clk  = \AES.r1.t3.t2.clk ;
    assign \AES.r1.t3.t2.s0.in  = \AES.r1.t3.t2.in ;
    assign \AES.r1.t3.t2.k0  = \AES.r1.t3.t2.s0.out ;
    always @ (  posedge \AES.r1.t3.t2.s0.clk )
    begin
        case ( \AES.r1.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t2.s4.clk  = \AES.r1.t3.t2.clk ;
    assign \AES.r1.t3.t2.s4.in  = \AES.r1.t3.t2.in ;
    assign \AES.r1.t3.t2.k1  = \AES.r1.t3.t2.s4.out ;
    always @ (  posedge \AES.r1.t3.t2.s4.clk )
    begin
        case ( \AES.r1.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t2.out  = { \AES.r1.t3.t2.k0 , \AES.r1.t3.t2.k0 , ( \AES.r1.t3.t2.k0  ^ \AES.r1.t3.t2.k1  ), \AES.r1.t3.t2.k1  };
    assign \AES.r1.t3.t3.clk  = \AES.r1.t3.clk ;
    assign \AES.r1.t3.t3.in  = \AES.r1.t3.b3 ;
    assign \AES.r1.t3.p3  = \AES.r1.t3.t3.out ;
    assign \AES.r1.t3.t3.s0.clk  = \AES.r1.t3.t3.clk ;
    assign \AES.r1.t3.t3.s0.in  = \AES.r1.t3.t3.in ;
    assign \AES.r1.t3.t3.k0  = \AES.r1.t3.t3.s0.out ;
    always @ (  posedge \AES.r1.t3.t3.s0.clk )
    begin
        case ( \AES.r1.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t3.s4.clk  = \AES.r1.t3.t3.clk ;
    assign \AES.r1.t3.t3.s4.in  = \AES.r1.t3.t3.in ;
    assign \AES.r1.t3.t3.k1  = \AES.r1.t3.t3.s4.out ;
    always @ (  posedge \AES.r1.t3.t3.s4.clk )
    begin
        case ( \AES.r1.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r1.t3.t3.out  = { \AES.r1.t3.t3.k0 , \AES.r1.t3.t3.k0 , ( \AES.r1.t3.t3.k0  ^ \AES.r1.t3.t3.k1  ), \AES.r1.t3.t3.k1  };
    assign \AES.r1.z0  = ( ( ( ( \AES.r1.p00  ^ \AES.r1.p11  ) ^ \AES.r1.p22  ) ^ \AES.r1.p33  ) ^ \AES.r1.k0  );
    assign \AES.r1.z1  = ( ( ( ( \AES.r1.p03  ^ \AES.r1.p10  ) ^ \AES.r1.p21  ) ^ \AES.r1.p32  ) ^ \AES.r1.k1  );
    assign \AES.r1.z2  = ( ( ( ( \AES.r1.p02  ^ \AES.r1.p13  ) ^ \AES.r1.p20  ) ^ \AES.r1.p31  ) ^ \AES.r1.k2  );
    assign \AES.r1.z3  = ( ( ( ( \AES.r1.p01  ^ \AES.r1.p12  ) ^ \AES.r1.p23  ) ^ \AES.r1.p30  ) ^ \AES.r1.k3  );
    always @ (  posedge \AES.r1.clk )
    begin
    end
    assign \AES.r2.clk  = \AES.clk ;
    assign \AES.r2.state_in  = \AES.s1 ;
    assign \AES.r2.key  = \AES.k1b ;
    assign \AES.s2  = \AES.r2.state_out ;
    assign \AES.r2.k0  = \AES.r2.key [127:96];
    assign \AES.r2.k1  = \AES.r2.key [95:64];
    assign \AES.r2.k2  = \AES.r2.key [63:32];
    assign \AES.r2.k3  = \AES.r2.key [31:0];
    assign \AES.r2.s0  = \AES.r2.state_in [127:96];
    assign \AES.r2.s1  = \AES.r2.state_in [95:64];
    assign \AES.r2.s2  = \AES.r2.state_in [63:32];
    assign \AES.r2.s3  = \AES.r2.state_in [31:0];
    assign \AES.r2.t0.clk  = \AES.r2.clk ;
    assign \AES.r2.t0.state  = \AES.r2.s0 ;
    assign \AES.r2.p00  = \AES.r2.t0.p0 ;
    assign \AES.r2.p01  = \AES.r2.t0.p1 ;
    assign \AES.r2.p02  = \AES.r2.t0.p2 ;
    assign \AES.r2.p03  = \AES.r2.t0.p3 ;
    assign \AES.r2.t0.p0  = { \AES.r2.t0.k0 [7:0], \AES.r2.t0.k0 [31:8] };
    assign \AES.r2.t0.p1  = { \AES.r2.t0.k1 [15:0], \AES.r2.t0.k1 [31:16] };
    assign \AES.r2.t0.p2  = { \AES.r2.t0.k2 [23:0], \AES.r2.t0.k2 [31:24] };
    assign \AES.r2.t0.b0  = \AES.r2.t0.state [31:24];
    assign \AES.r2.t0.b1  = \AES.r2.t0.state [23:16];
    assign \AES.r2.t0.b2  = \AES.r2.t0.state [15:8];
    assign \AES.r2.t0.b3  = \AES.r2.t0.state [7:0];
    assign \AES.r2.t0.t0.clk  = \AES.r2.t0.clk ;
    assign \AES.r2.t0.t0.in  = \AES.r2.t0.b0 ;
    assign \AES.r2.t0.k0  = \AES.r2.t0.t0.out ;
    assign \AES.r2.t0.t0.s0.clk  = \AES.r2.t0.t0.clk ;
    assign \AES.r2.t0.t0.s0.in  = \AES.r2.t0.t0.in ;
    assign \AES.r2.t0.t0.k0  = \AES.r2.t0.t0.s0.out ;
    always @ (  posedge \AES.r2.t0.t0.s0.clk )
    begin
        case ( \AES.r2.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t0.s4.clk  = \AES.r2.t0.t0.clk ;
    assign \AES.r2.t0.t0.s4.in  = \AES.r2.t0.t0.in ;
    assign \AES.r2.t0.t0.k1  = \AES.r2.t0.t0.s4.out ;
    always @ (  posedge \AES.r2.t0.t0.s4.clk )
    begin
        case ( \AES.r2.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t0.out  = { \AES.r2.t0.t0.k0 , \AES.r2.t0.t0.k0 , ( \AES.r2.t0.t0.k0  ^ \AES.r2.t0.t0.k1  ), \AES.r2.t0.t0.k1  };
    assign \AES.r2.t0.t1.clk  = \AES.r2.t0.clk ;
    assign \AES.r2.t0.t1.in  = \AES.r2.t0.b1 ;
    assign \AES.r2.t0.k1  = \AES.r2.t0.t1.out ;
    assign \AES.r2.t0.t1.s0.clk  = \AES.r2.t0.t1.clk ;
    assign \AES.r2.t0.t1.s0.in  = \AES.r2.t0.t1.in ;
    assign \AES.r2.t0.t1.k0  = \AES.r2.t0.t1.s0.out ;
    always @ (  posedge \AES.r2.t0.t1.s0.clk )
    begin
        case ( \AES.r2.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t1.s4.clk  = \AES.r2.t0.t1.clk ;
    assign \AES.r2.t0.t1.s4.in  = \AES.r2.t0.t1.in ;
    assign \AES.r2.t0.t1.k1  = \AES.r2.t0.t1.s4.out ;
    always @ (  posedge \AES.r2.t0.t1.s4.clk )
    begin
        case ( \AES.r2.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t1.out  = { \AES.r2.t0.t1.k0 , \AES.r2.t0.t1.k0 , ( \AES.r2.t0.t1.k0  ^ \AES.r2.t0.t1.k1  ), \AES.r2.t0.t1.k1  };
    assign \AES.r2.t0.t2.clk  = \AES.r2.t0.clk ;
    assign \AES.r2.t0.t2.in  = \AES.r2.t0.b2 ;
    assign \AES.r2.t0.k2  = \AES.r2.t0.t2.out ;
    assign \AES.r2.t0.t2.s0.clk  = \AES.r2.t0.t2.clk ;
    assign \AES.r2.t0.t2.s0.in  = \AES.r2.t0.t2.in ;
    assign \AES.r2.t0.t2.k0  = \AES.r2.t0.t2.s0.out ;
    always @ (  posedge \AES.r2.t0.t2.s0.clk )
    begin
        case ( \AES.r2.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t2.s4.clk  = \AES.r2.t0.t2.clk ;
    assign \AES.r2.t0.t2.s4.in  = \AES.r2.t0.t2.in ;
    assign \AES.r2.t0.t2.k1  = \AES.r2.t0.t2.s4.out ;
    always @ (  posedge \AES.r2.t0.t2.s4.clk )
    begin
        case ( \AES.r2.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t2.out  = { \AES.r2.t0.t2.k0 , \AES.r2.t0.t2.k0 , ( \AES.r2.t0.t2.k0  ^ \AES.r2.t0.t2.k1  ), \AES.r2.t0.t2.k1  };
    assign \AES.r2.t0.t3.clk  = \AES.r2.t0.clk ;
    assign \AES.r2.t0.t3.in  = \AES.r2.t0.b3 ;
    assign \AES.r2.t0.p3  = \AES.r2.t0.t3.out ;
    assign \AES.r2.t0.t3.s0.clk  = \AES.r2.t0.t3.clk ;
    assign \AES.r2.t0.t3.s0.in  = \AES.r2.t0.t3.in ;
    assign \AES.r2.t0.t3.k0  = \AES.r2.t0.t3.s0.out ;
    always @ (  posedge \AES.r2.t0.t3.s0.clk )
    begin
        case ( \AES.r2.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t3.s4.clk  = \AES.r2.t0.t3.clk ;
    assign \AES.r2.t0.t3.s4.in  = \AES.r2.t0.t3.in ;
    assign \AES.r2.t0.t3.k1  = \AES.r2.t0.t3.s4.out ;
    always @ (  posedge \AES.r2.t0.t3.s4.clk )
    begin
        case ( \AES.r2.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t0.t3.out  = { \AES.r2.t0.t3.k0 , \AES.r2.t0.t3.k0 , ( \AES.r2.t0.t3.k0  ^ \AES.r2.t0.t3.k1  ), \AES.r2.t0.t3.k1  };
    assign \AES.r2.t1.clk  = \AES.r2.clk ;
    assign \AES.r2.t1.state  = \AES.r2.s1 ;
    assign \AES.r2.p10  = \AES.r2.t1.p0 ;
    assign \AES.r2.p11  = \AES.r2.t1.p1 ;
    assign \AES.r2.p12  = \AES.r2.t1.p2 ;
    assign \AES.r2.p13  = \AES.r2.t1.p3 ;
    assign \AES.r2.t1.p0  = { \AES.r2.t1.k0 [7:0], \AES.r2.t1.k0 [31:8] };
    assign \AES.r2.t1.p1  = { \AES.r2.t1.k1 [15:0], \AES.r2.t1.k1 [31:16] };
    assign \AES.r2.t1.p2  = { \AES.r2.t1.k2 [23:0], \AES.r2.t1.k2 [31:24] };
    assign \AES.r2.t1.b0  = \AES.r2.t1.state [31:24];
    assign \AES.r2.t1.b1  = \AES.r2.t1.state [23:16];
    assign \AES.r2.t1.b2  = \AES.r2.t1.state [15:8];
    assign \AES.r2.t1.b3  = \AES.r2.t1.state [7:0];
    assign \AES.r2.t1.t0.clk  = \AES.r2.t1.clk ;
    assign \AES.r2.t1.t0.in  = \AES.r2.t1.b0 ;
    assign \AES.r2.t1.k0  = \AES.r2.t1.t0.out ;
    assign \AES.r2.t1.t0.s0.clk  = \AES.r2.t1.t0.clk ;
    assign \AES.r2.t1.t0.s0.in  = \AES.r2.t1.t0.in ;
    assign \AES.r2.t1.t0.k0  = \AES.r2.t1.t0.s0.out ;
    always @ (  posedge \AES.r2.t1.t0.s0.clk )
    begin
        case ( \AES.r2.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t0.s4.clk  = \AES.r2.t1.t0.clk ;
    assign \AES.r2.t1.t0.s4.in  = \AES.r2.t1.t0.in ;
    assign \AES.r2.t1.t0.k1  = \AES.r2.t1.t0.s4.out ;
    always @ (  posedge \AES.r2.t1.t0.s4.clk )
    begin
        case ( \AES.r2.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t0.out  = { \AES.r2.t1.t0.k0 , \AES.r2.t1.t0.k0 , ( \AES.r2.t1.t0.k0  ^ \AES.r2.t1.t0.k1  ), \AES.r2.t1.t0.k1  };
    assign \AES.r2.t1.t1.clk  = \AES.r2.t1.clk ;
    assign \AES.r2.t1.t1.in  = \AES.r2.t1.b1 ;
    assign \AES.r2.t1.k1  = \AES.r2.t1.t1.out ;
    assign \AES.r2.t1.t1.s0.clk  = \AES.r2.t1.t1.clk ;
    assign \AES.r2.t1.t1.s0.in  = \AES.r2.t1.t1.in ;
    assign \AES.r2.t1.t1.k0  = \AES.r2.t1.t1.s0.out ;
    always @ (  posedge \AES.r2.t1.t1.s0.clk )
    begin
        case ( \AES.r2.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t1.s4.clk  = \AES.r2.t1.t1.clk ;
    assign \AES.r2.t1.t1.s4.in  = \AES.r2.t1.t1.in ;
    assign \AES.r2.t1.t1.k1  = \AES.r2.t1.t1.s4.out ;
    always @ (  posedge \AES.r2.t1.t1.s4.clk )
    begin
        case ( \AES.r2.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t1.out  = { \AES.r2.t1.t1.k0 , \AES.r2.t1.t1.k0 , ( \AES.r2.t1.t1.k0  ^ \AES.r2.t1.t1.k1  ), \AES.r2.t1.t1.k1  };
    assign \AES.r2.t1.t2.clk  = \AES.r2.t1.clk ;
    assign \AES.r2.t1.t2.in  = \AES.r2.t1.b2 ;
    assign \AES.r2.t1.k2  = \AES.r2.t1.t2.out ;
    assign \AES.r2.t1.t2.s0.clk  = \AES.r2.t1.t2.clk ;
    assign \AES.r2.t1.t2.s0.in  = \AES.r2.t1.t2.in ;
    assign \AES.r2.t1.t2.k0  = \AES.r2.t1.t2.s0.out ;
    always @ (  posedge \AES.r2.t1.t2.s0.clk )
    begin
        case ( \AES.r2.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t2.s4.clk  = \AES.r2.t1.t2.clk ;
    assign \AES.r2.t1.t2.s4.in  = \AES.r2.t1.t2.in ;
    assign \AES.r2.t1.t2.k1  = \AES.r2.t1.t2.s4.out ;
    always @ (  posedge \AES.r2.t1.t2.s4.clk )
    begin
        case ( \AES.r2.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t2.out  = { \AES.r2.t1.t2.k0 , \AES.r2.t1.t2.k0 , ( \AES.r2.t1.t2.k0  ^ \AES.r2.t1.t2.k1  ), \AES.r2.t1.t2.k1  };
    assign \AES.r2.t1.t3.clk  = \AES.r2.t1.clk ;
    assign \AES.r2.t1.t3.in  = \AES.r2.t1.b3 ;
    assign \AES.r2.t1.p3  = \AES.r2.t1.t3.out ;
    assign \AES.r2.t1.t3.s0.clk  = \AES.r2.t1.t3.clk ;
    assign \AES.r2.t1.t3.s0.in  = \AES.r2.t1.t3.in ;
    assign \AES.r2.t1.t3.k0  = \AES.r2.t1.t3.s0.out ;
    always @ (  posedge \AES.r2.t1.t3.s0.clk )
    begin
        case ( \AES.r2.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t3.s4.clk  = \AES.r2.t1.t3.clk ;
    assign \AES.r2.t1.t3.s4.in  = \AES.r2.t1.t3.in ;
    assign \AES.r2.t1.t3.k1  = \AES.r2.t1.t3.s4.out ;
    always @ (  posedge \AES.r2.t1.t3.s4.clk )
    begin
        case ( \AES.r2.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t1.t3.out  = { \AES.r2.t1.t3.k0 , \AES.r2.t1.t3.k0 , ( \AES.r2.t1.t3.k0  ^ \AES.r2.t1.t3.k1  ), \AES.r2.t1.t3.k1  };
    assign \AES.r2.t2.clk  = \AES.r2.clk ;
    assign \AES.r2.t2.state  = \AES.r2.s2 ;
    assign \AES.r2.p20  = \AES.r2.t2.p0 ;
    assign \AES.r2.p21  = \AES.r2.t2.p1 ;
    assign \AES.r2.p22  = \AES.r2.t2.p2 ;
    assign \AES.r2.p23  = \AES.r2.t2.p3 ;
    assign \AES.r2.t2.p0  = { \AES.r2.t2.k0 [7:0], \AES.r2.t2.k0 [31:8] };
    assign \AES.r2.t2.p1  = { \AES.r2.t2.k1 [15:0], \AES.r2.t2.k1 [31:16] };
    assign \AES.r2.t2.p2  = { \AES.r2.t2.k2 [23:0], \AES.r2.t2.k2 [31:24] };
    assign \AES.r2.t2.b0  = \AES.r2.t2.state [31:24];
    assign \AES.r2.t2.b1  = \AES.r2.t2.state [23:16];
    assign \AES.r2.t2.b2  = \AES.r2.t2.state [15:8];
    assign \AES.r2.t2.b3  = \AES.r2.t2.state [7:0];
    assign \AES.r2.t2.t0.clk  = \AES.r2.t2.clk ;
    assign \AES.r2.t2.t0.in  = \AES.r2.t2.b0 ;
    assign \AES.r2.t2.k0  = \AES.r2.t2.t0.out ;
    assign \AES.r2.t2.t0.s0.clk  = \AES.r2.t2.t0.clk ;
    assign \AES.r2.t2.t0.s0.in  = \AES.r2.t2.t0.in ;
    assign \AES.r2.t2.t0.k0  = \AES.r2.t2.t0.s0.out ;
    always @ (  posedge \AES.r2.t2.t0.s0.clk )
    begin
        case ( \AES.r2.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t0.s4.clk  = \AES.r2.t2.t0.clk ;
    assign \AES.r2.t2.t0.s4.in  = \AES.r2.t2.t0.in ;
    assign \AES.r2.t2.t0.k1  = \AES.r2.t2.t0.s4.out ;
    always @ (  posedge \AES.r2.t2.t0.s4.clk )
    begin
        case ( \AES.r2.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t0.out  = { \AES.r2.t2.t0.k0 , \AES.r2.t2.t0.k0 , ( \AES.r2.t2.t0.k0  ^ \AES.r2.t2.t0.k1  ), \AES.r2.t2.t0.k1  };
    assign \AES.r2.t2.t1.clk  = \AES.r2.t2.clk ;
    assign \AES.r2.t2.t1.in  = \AES.r2.t2.b1 ;
    assign \AES.r2.t2.k1  = \AES.r2.t2.t1.out ;
    assign \AES.r2.t2.t1.s0.clk  = \AES.r2.t2.t1.clk ;
    assign \AES.r2.t2.t1.s0.in  = \AES.r2.t2.t1.in ;
    assign \AES.r2.t2.t1.k0  = \AES.r2.t2.t1.s0.out ;
    always @ (  posedge \AES.r2.t2.t1.s0.clk )
    begin
        case ( \AES.r2.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t1.s4.clk  = \AES.r2.t2.t1.clk ;
    assign \AES.r2.t2.t1.s4.in  = \AES.r2.t2.t1.in ;
    assign \AES.r2.t2.t1.k1  = \AES.r2.t2.t1.s4.out ;
    always @ (  posedge \AES.r2.t2.t1.s4.clk )
    begin
        case ( \AES.r2.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t1.out  = { \AES.r2.t2.t1.k0 , \AES.r2.t2.t1.k0 , ( \AES.r2.t2.t1.k0  ^ \AES.r2.t2.t1.k1  ), \AES.r2.t2.t1.k1  };
    assign \AES.r2.t2.t2.clk  = \AES.r2.t2.clk ;
    assign \AES.r2.t2.t2.in  = \AES.r2.t2.b2 ;
    assign \AES.r2.t2.k2  = \AES.r2.t2.t2.out ;
    assign \AES.r2.t2.t2.s0.clk  = \AES.r2.t2.t2.clk ;
    assign \AES.r2.t2.t2.s0.in  = \AES.r2.t2.t2.in ;
    assign \AES.r2.t2.t2.k0  = \AES.r2.t2.t2.s0.out ;
    always @ (  posedge \AES.r2.t2.t2.s0.clk )
    begin
        case ( \AES.r2.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t2.s4.clk  = \AES.r2.t2.t2.clk ;
    assign \AES.r2.t2.t2.s4.in  = \AES.r2.t2.t2.in ;
    assign \AES.r2.t2.t2.k1  = \AES.r2.t2.t2.s4.out ;
    always @ (  posedge \AES.r2.t2.t2.s4.clk )
    begin
        case ( \AES.r2.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t2.out  = { \AES.r2.t2.t2.k0 , \AES.r2.t2.t2.k0 , ( \AES.r2.t2.t2.k0  ^ \AES.r2.t2.t2.k1  ), \AES.r2.t2.t2.k1  };
    assign \AES.r2.t2.t3.clk  = \AES.r2.t2.clk ;
    assign \AES.r2.t2.t3.in  = \AES.r2.t2.b3 ;
    assign \AES.r2.t2.p3  = \AES.r2.t2.t3.out ;
    assign \AES.r2.t2.t3.s0.clk  = \AES.r2.t2.t3.clk ;
    assign \AES.r2.t2.t3.s0.in  = \AES.r2.t2.t3.in ;
    assign \AES.r2.t2.t3.k0  = \AES.r2.t2.t3.s0.out ;
    always @ (  posedge \AES.r2.t2.t3.s0.clk )
    begin
        case ( \AES.r2.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t3.s4.clk  = \AES.r2.t2.t3.clk ;
    assign \AES.r2.t2.t3.s4.in  = \AES.r2.t2.t3.in ;
    assign \AES.r2.t2.t3.k1  = \AES.r2.t2.t3.s4.out ;
    always @ (  posedge \AES.r2.t2.t3.s4.clk )
    begin
        case ( \AES.r2.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t2.t3.out  = { \AES.r2.t2.t3.k0 , \AES.r2.t2.t3.k0 , ( \AES.r2.t2.t3.k0  ^ \AES.r2.t2.t3.k1  ), \AES.r2.t2.t3.k1  };
    assign \AES.r2.t3.clk  = \AES.r2.clk ;
    assign \AES.r2.t3.state  = \AES.r2.s3 ;
    assign \AES.r2.p30  = \AES.r2.t3.p0 ;
    assign \AES.r2.p31  = \AES.r2.t3.p1 ;
    assign \AES.r2.p32  = \AES.r2.t3.p2 ;
    assign \AES.r2.p33  = \AES.r2.t3.p3 ;
    assign \AES.r2.t3.p0  = { \AES.r2.t3.k0 [7:0], \AES.r2.t3.k0 [31:8] };
    assign \AES.r2.t3.p1  = { \AES.r2.t3.k1 [15:0], \AES.r2.t3.k1 [31:16] };
    assign \AES.r2.t3.p2  = { \AES.r2.t3.k2 [23:0], \AES.r2.t3.k2 [31:24] };
    assign \AES.r2.t3.b0  = \AES.r2.t3.state [31:24];
    assign \AES.r2.t3.b1  = \AES.r2.t3.state [23:16];
    assign \AES.r2.t3.b2  = \AES.r2.t3.state [15:8];
    assign \AES.r2.t3.b3  = \AES.r2.t3.state [7:0];
    assign \AES.r2.t3.t0.clk  = \AES.r2.t3.clk ;
    assign \AES.r2.t3.t0.in  = \AES.r2.t3.b0 ;
    assign \AES.r2.t3.k0  = \AES.r2.t3.t0.out ;
    assign \AES.r2.t3.t0.s0.clk  = \AES.r2.t3.t0.clk ;
    assign \AES.r2.t3.t0.s0.in  = \AES.r2.t3.t0.in ;
    assign \AES.r2.t3.t0.k0  = \AES.r2.t3.t0.s0.out ;
    always @ (  posedge \AES.r2.t3.t0.s0.clk )
    begin
        case ( \AES.r2.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t0.s4.clk  = \AES.r2.t3.t0.clk ;
    assign \AES.r2.t3.t0.s4.in  = \AES.r2.t3.t0.in ;
    assign \AES.r2.t3.t0.k1  = \AES.r2.t3.t0.s4.out ;
    always @ (  posedge \AES.r2.t3.t0.s4.clk )
    begin
        case ( \AES.r2.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t0.out  = { \AES.r2.t3.t0.k0 , \AES.r2.t3.t0.k0 , ( \AES.r2.t3.t0.k0  ^ \AES.r2.t3.t0.k1  ), \AES.r2.t3.t0.k1  };
    assign \AES.r2.t3.t1.clk  = \AES.r2.t3.clk ;
    assign \AES.r2.t3.t1.in  = \AES.r2.t3.b1 ;
    assign \AES.r2.t3.k1  = \AES.r2.t3.t1.out ;
    assign \AES.r2.t3.t1.s0.clk  = \AES.r2.t3.t1.clk ;
    assign \AES.r2.t3.t1.s0.in  = \AES.r2.t3.t1.in ;
    assign \AES.r2.t3.t1.k0  = \AES.r2.t3.t1.s0.out ;
    always @ (  posedge \AES.r2.t3.t1.s0.clk )
    begin
        case ( \AES.r2.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t1.s4.clk  = \AES.r2.t3.t1.clk ;
    assign \AES.r2.t3.t1.s4.in  = \AES.r2.t3.t1.in ;
    assign \AES.r2.t3.t1.k1  = \AES.r2.t3.t1.s4.out ;
    always @ (  posedge \AES.r2.t3.t1.s4.clk )
    begin
        case ( \AES.r2.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t1.out  = { \AES.r2.t3.t1.k0 , \AES.r2.t3.t1.k0 , ( \AES.r2.t3.t1.k0  ^ \AES.r2.t3.t1.k1  ), \AES.r2.t3.t1.k1  };
    assign \AES.r2.t3.t2.clk  = \AES.r2.t3.clk ;
    assign \AES.r2.t3.t2.in  = \AES.r2.t3.b2 ;
    assign \AES.r2.t3.k2  = \AES.r2.t3.t2.out ;
    assign \AES.r2.t3.t2.s0.clk  = \AES.r2.t3.t2.clk ;
    assign \AES.r2.t3.t2.s0.in  = \AES.r2.t3.t2.in ;
    assign \AES.r2.t3.t2.k0  = \AES.r2.t3.t2.s0.out ;
    always @ (  posedge \AES.r2.t3.t2.s0.clk )
    begin
        case ( \AES.r2.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t2.s4.clk  = \AES.r2.t3.t2.clk ;
    assign \AES.r2.t3.t2.s4.in  = \AES.r2.t3.t2.in ;
    assign \AES.r2.t3.t2.k1  = \AES.r2.t3.t2.s4.out ;
    always @ (  posedge \AES.r2.t3.t2.s4.clk )
    begin
        case ( \AES.r2.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t2.out  = { \AES.r2.t3.t2.k0 , \AES.r2.t3.t2.k0 , ( \AES.r2.t3.t2.k0  ^ \AES.r2.t3.t2.k1  ), \AES.r2.t3.t2.k1  };
    assign \AES.r2.t3.t3.clk  = \AES.r2.t3.clk ;
    assign \AES.r2.t3.t3.in  = \AES.r2.t3.b3 ;
    assign \AES.r2.t3.p3  = \AES.r2.t3.t3.out ;
    assign \AES.r2.t3.t3.s0.clk  = \AES.r2.t3.t3.clk ;
    assign \AES.r2.t3.t3.s0.in  = \AES.r2.t3.t3.in ;
    assign \AES.r2.t3.t3.k0  = \AES.r2.t3.t3.s0.out ;
    always @ (  posedge \AES.r2.t3.t3.s0.clk )
    begin
        case ( \AES.r2.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t3.s4.clk  = \AES.r2.t3.t3.clk ;
    assign \AES.r2.t3.t3.s4.in  = \AES.r2.t3.t3.in ;
    assign \AES.r2.t3.t3.k1  = \AES.r2.t3.t3.s4.out ;
    always @ (  posedge \AES.r2.t3.t3.s4.clk )
    begin
        case ( \AES.r2.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r2.t3.t3.out  = { \AES.r2.t3.t3.k0 , \AES.r2.t3.t3.k0 , ( \AES.r2.t3.t3.k0  ^ \AES.r2.t3.t3.k1  ), \AES.r2.t3.t3.k1  };
    assign \AES.r2.z0  = ( ( ( ( \AES.r2.p00  ^ \AES.r2.p11  ) ^ \AES.r2.p22  ) ^ \AES.r2.p33  ) ^ \AES.r2.k0  );
    assign \AES.r2.z1  = ( ( ( ( \AES.r2.p03  ^ \AES.r2.p10  ) ^ \AES.r2.p21  ) ^ \AES.r2.p32  ) ^ \AES.r2.k1  );
    assign \AES.r2.z2  = ( ( ( ( \AES.r2.p02  ^ \AES.r2.p13  ) ^ \AES.r2.p20  ) ^ \AES.r2.p31  ) ^ \AES.r2.k2  );
    assign \AES.r2.z3  = ( ( ( ( \AES.r2.p01  ^ \AES.r2.p12  ) ^ \AES.r2.p23  ) ^ \AES.r2.p30  ) ^ \AES.r2.k3  );
    always @ (  posedge \AES.r2.clk )
    begin
    end
    assign \AES.r3.clk  = \AES.clk ;
    assign \AES.r3.state_in  = \AES.s2 ;
    assign \AES.r3.key  = \AES.k2b ;
    assign \AES.s3  = \AES.r3.state_out ;
    assign \AES.r3.k0  = \AES.r3.key [127:96];
    assign \AES.r3.k1  = \AES.r3.key [95:64];
    assign \AES.r3.k2  = \AES.r3.key [63:32];
    assign \AES.r3.k3  = \AES.r3.key [31:0];
    assign \AES.r3.s0  = \AES.r3.state_in [127:96];
    assign \AES.r3.s1  = \AES.r3.state_in [95:64];
    assign \AES.r3.s2  = \AES.r3.state_in [63:32];
    assign \AES.r3.s3  = \AES.r3.state_in [31:0];
    assign \AES.r3.t0.clk  = \AES.r3.clk ;
    assign \AES.r3.t0.state  = \AES.r3.s0 ;
    assign \AES.r3.p00  = \AES.r3.t0.p0 ;
    assign \AES.r3.p01  = \AES.r3.t0.p1 ;
    assign \AES.r3.p02  = \AES.r3.t0.p2 ;
    assign \AES.r3.p03  = \AES.r3.t0.p3 ;
    assign \AES.r3.t0.p0  = { \AES.r3.t0.k0 [7:0], \AES.r3.t0.k0 [31:8] };
    assign \AES.r3.t0.p1  = { \AES.r3.t0.k1 [15:0], \AES.r3.t0.k1 [31:16] };
    assign \AES.r3.t0.p2  = { \AES.r3.t0.k2 [23:0], \AES.r3.t0.k2 [31:24] };
    assign \AES.r3.t0.b0  = \AES.r3.t0.state [31:24];
    assign \AES.r3.t0.b1  = \AES.r3.t0.state [23:16];
    assign \AES.r3.t0.b2  = \AES.r3.t0.state [15:8];
    assign \AES.r3.t0.b3  = \AES.r3.t0.state [7:0];
    assign \AES.r3.t0.t0.clk  = \AES.r3.t0.clk ;
    assign \AES.r3.t0.t0.in  = \AES.r3.t0.b0 ;
    assign \AES.r3.t0.k0  = \AES.r3.t0.t0.out ;
    assign \AES.r3.t0.t0.s0.clk  = \AES.r3.t0.t0.clk ;
    assign \AES.r3.t0.t0.s0.in  = \AES.r3.t0.t0.in ;
    assign \AES.r3.t0.t0.k0  = \AES.r3.t0.t0.s0.out ;
    always @ (  posedge \AES.r3.t0.t0.s0.clk )
    begin
        case ( \AES.r3.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t0.s4.clk  = \AES.r3.t0.t0.clk ;
    assign \AES.r3.t0.t0.s4.in  = \AES.r3.t0.t0.in ;
    assign \AES.r3.t0.t0.k1  = \AES.r3.t0.t0.s4.out ;
    always @ (  posedge \AES.r3.t0.t0.s4.clk )
    begin
        case ( \AES.r3.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t0.out  = { \AES.r3.t0.t0.k0 , \AES.r3.t0.t0.k0 , ( \AES.r3.t0.t0.k0  ^ \AES.r3.t0.t0.k1  ), \AES.r3.t0.t0.k1  };
    assign \AES.r3.t0.t1.clk  = \AES.r3.t0.clk ;
    assign \AES.r3.t0.t1.in  = \AES.r3.t0.b1 ;
    assign \AES.r3.t0.k1  = \AES.r3.t0.t1.out ;
    assign \AES.r3.t0.t1.s0.clk  = \AES.r3.t0.t1.clk ;
    assign \AES.r3.t0.t1.s0.in  = \AES.r3.t0.t1.in ;
    assign \AES.r3.t0.t1.k0  = \AES.r3.t0.t1.s0.out ;
    always @ (  posedge \AES.r3.t0.t1.s0.clk )
    begin
        case ( \AES.r3.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t1.s4.clk  = \AES.r3.t0.t1.clk ;
    assign \AES.r3.t0.t1.s4.in  = \AES.r3.t0.t1.in ;
    assign \AES.r3.t0.t1.k1  = \AES.r3.t0.t1.s4.out ;
    always @ (  posedge \AES.r3.t0.t1.s4.clk )
    begin
        case ( \AES.r3.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t1.out  = { \AES.r3.t0.t1.k0 , \AES.r3.t0.t1.k0 , ( \AES.r3.t0.t1.k0  ^ \AES.r3.t0.t1.k1  ), \AES.r3.t0.t1.k1  };
    assign \AES.r3.t0.t2.clk  = \AES.r3.t0.clk ;
    assign \AES.r3.t0.t2.in  = \AES.r3.t0.b2 ;
    assign \AES.r3.t0.k2  = \AES.r3.t0.t2.out ;
    assign \AES.r3.t0.t2.s0.clk  = \AES.r3.t0.t2.clk ;
    assign \AES.r3.t0.t2.s0.in  = \AES.r3.t0.t2.in ;
    assign \AES.r3.t0.t2.k0  = \AES.r3.t0.t2.s0.out ;
    always @ (  posedge \AES.r3.t0.t2.s0.clk )
    begin
        case ( \AES.r3.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t2.s4.clk  = \AES.r3.t0.t2.clk ;
    assign \AES.r3.t0.t2.s4.in  = \AES.r3.t0.t2.in ;
    assign \AES.r3.t0.t2.k1  = \AES.r3.t0.t2.s4.out ;
    always @ (  posedge \AES.r3.t0.t2.s4.clk )
    begin
        case ( \AES.r3.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t2.out  = { \AES.r3.t0.t2.k0 , \AES.r3.t0.t2.k0 , ( \AES.r3.t0.t2.k0  ^ \AES.r3.t0.t2.k1  ), \AES.r3.t0.t2.k1  };
    assign \AES.r3.t0.t3.clk  = \AES.r3.t0.clk ;
    assign \AES.r3.t0.t3.in  = \AES.r3.t0.b3 ;
    assign \AES.r3.t0.p3  = \AES.r3.t0.t3.out ;
    assign \AES.r3.t0.t3.s0.clk  = \AES.r3.t0.t3.clk ;
    assign \AES.r3.t0.t3.s0.in  = \AES.r3.t0.t3.in ;
    assign \AES.r3.t0.t3.k0  = \AES.r3.t0.t3.s0.out ;
    always @ (  posedge \AES.r3.t0.t3.s0.clk )
    begin
        case ( \AES.r3.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t3.s4.clk  = \AES.r3.t0.t3.clk ;
    assign \AES.r3.t0.t3.s4.in  = \AES.r3.t0.t3.in ;
    assign \AES.r3.t0.t3.k1  = \AES.r3.t0.t3.s4.out ;
    always @ (  posedge \AES.r3.t0.t3.s4.clk )
    begin
        case ( \AES.r3.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t0.t3.out  = { \AES.r3.t0.t3.k0 , \AES.r3.t0.t3.k0 , ( \AES.r3.t0.t3.k0  ^ \AES.r3.t0.t3.k1  ), \AES.r3.t0.t3.k1  };
    assign \AES.r3.t1.clk  = \AES.r3.clk ;
    assign \AES.r3.t1.state  = \AES.r3.s1 ;
    assign \AES.r3.p10  = \AES.r3.t1.p0 ;
    assign \AES.r3.p11  = \AES.r3.t1.p1 ;
    assign \AES.r3.p12  = \AES.r3.t1.p2 ;
    assign \AES.r3.p13  = \AES.r3.t1.p3 ;
    assign \AES.r3.t1.p0  = { \AES.r3.t1.k0 [7:0], \AES.r3.t1.k0 [31:8] };
    assign \AES.r3.t1.p1  = { \AES.r3.t1.k1 [15:0], \AES.r3.t1.k1 [31:16] };
    assign \AES.r3.t1.p2  = { \AES.r3.t1.k2 [23:0], \AES.r3.t1.k2 [31:24] };
    assign \AES.r3.t1.b0  = \AES.r3.t1.state [31:24];
    assign \AES.r3.t1.b1  = \AES.r3.t1.state [23:16];
    assign \AES.r3.t1.b2  = \AES.r3.t1.state [15:8];
    assign \AES.r3.t1.b3  = \AES.r3.t1.state [7:0];
    assign \AES.r3.t1.t0.clk  = \AES.r3.t1.clk ;
    assign \AES.r3.t1.t0.in  = \AES.r3.t1.b0 ;
    assign \AES.r3.t1.k0  = \AES.r3.t1.t0.out ;
    assign \AES.r3.t1.t0.s0.clk  = \AES.r3.t1.t0.clk ;
    assign \AES.r3.t1.t0.s0.in  = \AES.r3.t1.t0.in ;
    assign \AES.r3.t1.t0.k0  = \AES.r3.t1.t0.s0.out ;
    always @ (  posedge \AES.r3.t1.t0.s0.clk )
    begin
        case ( \AES.r3.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t0.s4.clk  = \AES.r3.t1.t0.clk ;
    assign \AES.r3.t1.t0.s4.in  = \AES.r3.t1.t0.in ;
    assign \AES.r3.t1.t0.k1  = \AES.r3.t1.t0.s4.out ;
    always @ (  posedge \AES.r3.t1.t0.s4.clk )
    begin
        case ( \AES.r3.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t0.out  = { \AES.r3.t1.t0.k0 , \AES.r3.t1.t0.k0 , ( \AES.r3.t1.t0.k0  ^ \AES.r3.t1.t0.k1  ), \AES.r3.t1.t0.k1  };
    assign \AES.r3.t1.t1.clk  = \AES.r3.t1.clk ;
    assign \AES.r3.t1.t1.in  = \AES.r3.t1.b1 ;
    assign \AES.r3.t1.k1  = \AES.r3.t1.t1.out ;
    assign \AES.r3.t1.t1.s0.clk  = \AES.r3.t1.t1.clk ;
    assign \AES.r3.t1.t1.s0.in  = \AES.r3.t1.t1.in ;
    assign \AES.r3.t1.t1.k0  = \AES.r3.t1.t1.s0.out ;
    always @ (  posedge \AES.r3.t1.t1.s0.clk )
    begin
        case ( \AES.r3.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t1.s4.clk  = \AES.r3.t1.t1.clk ;
    assign \AES.r3.t1.t1.s4.in  = \AES.r3.t1.t1.in ;
    assign \AES.r3.t1.t1.k1  = \AES.r3.t1.t1.s4.out ;
    always @ (  posedge \AES.r3.t1.t1.s4.clk )
    begin
        case ( \AES.r3.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t1.out  = { \AES.r3.t1.t1.k0 , \AES.r3.t1.t1.k0 , ( \AES.r3.t1.t1.k0  ^ \AES.r3.t1.t1.k1  ), \AES.r3.t1.t1.k1  };
    assign \AES.r3.t1.t2.clk  = \AES.r3.t1.clk ;
    assign \AES.r3.t1.t2.in  = \AES.r3.t1.b2 ;
    assign \AES.r3.t1.k2  = \AES.r3.t1.t2.out ;
    assign \AES.r3.t1.t2.s0.clk  = \AES.r3.t1.t2.clk ;
    assign \AES.r3.t1.t2.s0.in  = \AES.r3.t1.t2.in ;
    assign \AES.r3.t1.t2.k0  = \AES.r3.t1.t2.s0.out ;
    always @ (  posedge \AES.r3.t1.t2.s0.clk )
    begin
        case ( \AES.r3.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t2.s4.clk  = \AES.r3.t1.t2.clk ;
    assign \AES.r3.t1.t2.s4.in  = \AES.r3.t1.t2.in ;
    assign \AES.r3.t1.t2.k1  = \AES.r3.t1.t2.s4.out ;
    always @ (  posedge \AES.r3.t1.t2.s4.clk )
    begin
        case ( \AES.r3.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t2.out  = { \AES.r3.t1.t2.k0 , \AES.r3.t1.t2.k0 , ( \AES.r3.t1.t2.k0  ^ \AES.r3.t1.t2.k1  ), \AES.r3.t1.t2.k1  };
    assign \AES.r3.t1.t3.clk  = \AES.r3.t1.clk ;
    assign \AES.r3.t1.t3.in  = \AES.r3.t1.b3 ;
    assign \AES.r3.t1.p3  = \AES.r3.t1.t3.out ;
    assign \AES.r3.t1.t3.s0.clk  = \AES.r3.t1.t3.clk ;
    assign \AES.r3.t1.t3.s0.in  = \AES.r3.t1.t3.in ;
    assign \AES.r3.t1.t3.k0  = \AES.r3.t1.t3.s0.out ;
    always @ (  posedge \AES.r3.t1.t3.s0.clk )
    begin
        case ( \AES.r3.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t3.s4.clk  = \AES.r3.t1.t3.clk ;
    assign \AES.r3.t1.t3.s4.in  = \AES.r3.t1.t3.in ;
    assign \AES.r3.t1.t3.k1  = \AES.r3.t1.t3.s4.out ;
    always @ (  posedge \AES.r3.t1.t3.s4.clk )
    begin
        case ( \AES.r3.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t1.t3.out  = { \AES.r3.t1.t3.k0 , \AES.r3.t1.t3.k0 , ( \AES.r3.t1.t3.k0  ^ \AES.r3.t1.t3.k1  ), \AES.r3.t1.t3.k1  };
    assign \AES.r3.t2.clk  = \AES.r3.clk ;
    assign \AES.r3.t2.state  = \AES.r3.s2 ;
    assign \AES.r3.p20  = \AES.r3.t2.p0 ;
    assign \AES.r3.p21  = \AES.r3.t2.p1 ;
    assign \AES.r3.p22  = \AES.r3.t2.p2 ;
    assign \AES.r3.p23  = \AES.r3.t2.p3 ;
    assign \AES.r3.t2.p0  = { \AES.r3.t2.k0 [7:0], \AES.r3.t2.k0 [31:8] };
    assign \AES.r3.t2.p1  = { \AES.r3.t2.k1 [15:0], \AES.r3.t2.k1 [31:16] };
    assign \AES.r3.t2.p2  = { \AES.r3.t2.k2 [23:0], \AES.r3.t2.k2 [31:24] };
    assign \AES.r3.t2.b0  = \AES.r3.t2.state [31:24];
    assign \AES.r3.t2.b1  = \AES.r3.t2.state [23:16];
    assign \AES.r3.t2.b2  = \AES.r3.t2.state [15:8];
    assign \AES.r3.t2.b3  = \AES.r3.t2.state [7:0];
    assign \AES.r3.t2.t0.clk  = \AES.r3.t2.clk ;
    assign \AES.r3.t2.t0.in  = \AES.r3.t2.b0 ;
    assign \AES.r3.t2.k0  = \AES.r3.t2.t0.out ;
    assign \AES.r3.t2.t0.s0.clk  = \AES.r3.t2.t0.clk ;
    assign \AES.r3.t2.t0.s0.in  = \AES.r3.t2.t0.in ;
    assign \AES.r3.t2.t0.k0  = \AES.r3.t2.t0.s0.out ;
    always @ (  posedge \AES.r3.t2.t0.s0.clk )
    begin
        case ( \AES.r3.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t0.s4.clk  = \AES.r3.t2.t0.clk ;
    assign \AES.r3.t2.t0.s4.in  = \AES.r3.t2.t0.in ;
    assign \AES.r3.t2.t0.k1  = \AES.r3.t2.t0.s4.out ;
    always @ (  posedge \AES.r3.t2.t0.s4.clk )
    begin
        case ( \AES.r3.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t0.out  = { \AES.r3.t2.t0.k0 , \AES.r3.t2.t0.k0 , ( \AES.r3.t2.t0.k0  ^ \AES.r3.t2.t0.k1  ), \AES.r3.t2.t0.k1  };
    assign \AES.r3.t2.t1.clk  = \AES.r3.t2.clk ;
    assign \AES.r3.t2.t1.in  = \AES.r3.t2.b1 ;
    assign \AES.r3.t2.k1  = \AES.r3.t2.t1.out ;
    assign \AES.r3.t2.t1.s0.clk  = \AES.r3.t2.t1.clk ;
    assign \AES.r3.t2.t1.s0.in  = \AES.r3.t2.t1.in ;
    assign \AES.r3.t2.t1.k0  = \AES.r3.t2.t1.s0.out ;
    always @ (  posedge \AES.r3.t2.t1.s0.clk )
    begin
        case ( \AES.r3.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t1.s4.clk  = \AES.r3.t2.t1.clk ;
    assign \AES.r3.t2.t1.s4.in  = \AES.r3.t2.t1.in ;
    assign \AES.r3.t2.t1.k1  = \AES.r3.t2.t1.s4.out ;
    always @ (  posedge \AES.r3.t2.t1.s4.clk )
    begin
        case ( \AES.r3.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t1.out  = { \AES.r3.t2.t1.k0 , \AES.r3.t2.t1.k0 , ( \AES.r3.t2.t1.k0  ^ \AES.r3.t2.t1.k1  ), \AES.r3.t2.t1.k1  };
    assign \AES.r3.t2.t2.clk  = \AES.r3.t2.clk ;
    assign \AES.r3.t2.t2.in  = \AES.r3.t2.b2 ;
    assign \AES.r3.t2.k2  = \AES.r3.t2.t2.out ;
    assign \AES.r3.t2.t2.s0.clk  = \AES.r3.t2.t2.clk ;
    assign \AES.r3.t2.t2.s0.in  = \AES.r3.t2.t2.in ;
    assign \AES.r3.t2.t2.k0  = \AES.r3.t2.t2.s0.out ;
    always @ (  posedge \AES.r3.t2.t2.s0.clk )
    begin
        case ( \AES.r3.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t2.s4.clk  = \AES.r3.t2.t2.clk ;
    assign \AES.r3.t2.t2.s4.in  = \AES.r3.t2.t2.in ;
    assign \AES.r3.t2.t2.k1  = \AES.r3.t2.t2.s4.out ;
    always @ (  posedge \AES.r3.t2.t2.s4.clk )
    begin
        case ( \AES.r3.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t2.out  = { \AES.r3.t2.t2.k0 , \AES.r3.t2.t2.k0 , ( \AES.r3.t2.t2.k0  ^ \AES.r3.t2.t2.k1  ), \AES.r3.t2.t2.k1  };
    assign \AES.r3.t2.t3.clk  = \AES.r3.t2.clk ;
    assign \AES.r3.t2.t3.in  = \AES.r3.t2.b3 ;
    assign \AES.r3.t2.p3  = \AES.r3.t2.t3.out ;
    assign \AES.r3.t2.t3.s0.clk  = \AES.r3.t2.t3.clk ;
    assign \AES.r3.t2.t3.s0.in  = \AES.r3.t2.t3.in ;
    assign \AES.r3.t2.t3.k0  = \AES.r3.t2.t3.s0.out ;
    always @ (  posedge \AES.r3.t2.t3.s0.clk )
    begin
        case ( \AES.r3.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t3.s4.clk  = \AES.r3.t2.t3.clk ;
    assign \AES.r3.t2.t3.s4.in  = \AES.r3.t2.t3.in ;
    assign \AES.r3.t2.t3.k1  = \AES.r3.t2.t3.s4.out ;
    always @ (  posedge \AES.r3.t2.t3.s4.clk )
    begin
        case ( \AES.r3.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t2.t3.out  = { \AES.r3.t2.t3.k0 , \AES.r3.t2.t3.k0 , ( \AES.r3.t2.t3.k0  ^ \AES.r3.t2.t3.k1  ), \AES.r3.t2.t3.k1  };
    assign \AES.r3.t3.clk  = \AES.r3.clk ;
    assign \AES.r3.t3.state  = \AES.r3.s3 ;
    assign \AES.r3.p30  = \AES.r3.t3.p0 ;
    assign \AES.r3.p31  = \AES.r3.t3.p1 ;
    assign \AES.r3.p32  = \AES.r3.t3.p2 ;
    assign \AES.r3.p33  = \AES.r3.t3.p3 ;
    assign \AES.r3.t3.p0  = { \AES.r3.t3.k0 [7:0], \AES.r3.t3.k0 [31:8] };
    assign \AES.r3.t3.p1  = { \AES.r3.t3.k1 [15:0], \AES.r3.t3.k1 [31:16] };
    assign \AES.r3.t3.p2  = { \AES.r3.t3.k2 [23:0], \AES.r3.t3.k2 [31:24] };
    assign \AES.r3.t3.b0  = \AES.r3.t3.state [31:24];
    assign \AES.r3.t3.b1  = \AES.r3.t3.state [23:16];
    assign \AES.r3.t3.b2  = \AES.r3.t3.state [15:8];
    assign \AES.r3.t3.b3  = \AES.r3.t3.state [7:0];
    assign \AES.r3.t3.t0.clk  = \AES.r3.t3.clk ;
    assign \AES.r3.t3.t0.in  = \AES.r3.t3.b0 ;
    assign \AES.r3.t3.k0  = \AES.r3.t3.t0.out ;
    assign \AES.r3.t3.t0.s0.clk  = \AES.r3.t3.t0.clk ;
    assign \AES.r3.t3.t0.s0.in  = \AES.r3.t3.t0.in ;
    assign \AES.r3.t3.t0.k0  = \AES.r3.t3.t0.s0.out ;
    always @ (  posedge \AES.r3.t3.t0.s0.clk )
    begin
        case ( \AES.r3.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t0.s4.clk  = \AES.r3.t3.t0.clk ;
    assign \AES.r3.t3.t0.s4.in  = \AES.r3.t3.t0.in ;
    assign \AES.r3.t3.t0.k1  = \AES.r3.t3.t0.s4.out ;
    always @ (  posedge \AES.r3.t3.t0.s4.clk )
    begin
        case ( \AES.r3.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t0.out  = { \AES.r3.t3.t0.k0 , \AES.r3.t3.t0.k0 , ( \AES.r3.t3.t0.k0  ^ \AES.r3.t3.t0.k1  ), \AES.r3.t3.t0.k1  };
    assign \AES.r3.t3.t1.clk  = \AES.r3.t3.clk ;
    assign \AES.r3.t3.t1.in  = \AES.r3.t3.b1 ;
    assign \AES.r3.t3.k1  = \AES.r3.t3.t1.out ;
    assign \AES.r3.t3.t1.s0.clk  = \AES.r3.t3.t1.clk ;
    assign \AES.r3.t3.t1.s0.in  = \AES.r3.t3.t1.in ;
    assign \AES.r3.t3.t1.k0  = \AES.r3.t3.t1.s0.out ;
    always @ (  posedge \AES.r3.t3.t1.s0.clk )
    begin
        case ( \AES.r3.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t1.s4.clk  = \AES.r3.t3.t1.clk ;
    assign \AES.r3.t3.t1.s4.in  = \AES.r3.t3.t1.in ;
    assign \AES.r3.t3.t1.k1  = \AES.r3.t3.t1.s4.out ;
    always @ (  posedge \AES.r3.t3.t1.s4.clk )
    begin
        case ( \AES.r3.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t1.out  = { \AES.r3.t3.t1.k0 , \AES.r3.t3.t1.k0 , ( \AES.r3.t3.t1.k0  ^ \AES.r3.t3.t1.k1  ), \AES.r3.t3.t1.k1  };
    assign \AES.r3.t3.t2.clk  = \AES.r3.t3.clk ;
    assign \AES.r3.t3.t2.in  = \AES.r3.t3.b2 ;
    assign \AES.r3.t3.k2  = \AES.r3.t3.t2.out ;
    assign \AES.r3.t3.t2.s0.clk  = \AES.r3.t3.t2.clk ;
    assign \AES.r3.t3.t2.s0.in  = \AES.r3.t3.t2.in ;
    assign \AES.r3.t3.t2.k0  = \AES.r3.t3.t2.s0.out ;
    always @ (  posedge \AES.r3.t3.t2.s0.clk )
    begin
        case ( \AES.r3.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t2.s4.clk  = \AES.r3.t3.t2.clk ;
    assign \AES.r3.t3.t2.s4.in  = \AES.r3.t3.t2.in ;
    assign \AES.r3.t3.t2.k1  = \AES.r3.t3.t2.s4.out ;
    always @ (  posedge \AES.r3.t3.t2.s4.clk )
    begin
        case ( \AES.r3.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t2.out  = { \AES.r3.t3.t2.k0 , \AES.r3.t3.t2.k0 , ( \AES.r3.t3.t2.k0  ^ \AES.r3.t3.t2.k1  ), \AES.r3.t3.t2.k1  };
    assign \AES.r3.t3.t3.clk  = \AES.r3.t3.clk ;
    assign \AES.r3.t3.t3.in  = \AES.r3.t3.b3 ;
    assign \AES.r3.t3.p3  = \AES.r3.t3.t3.out ;
    assign \AES.r3.t3.t3.s0.clk  = \AES.r3.t3.t3.clk ;
    assign \AES.r3.t3.t3.s0.in  = \AES.r3.t3.t3.in ;
    assign \AES.r3.t3.t3.k0  = \AES.r3.t3.t3.s0.out ;
    always @ (  posedge \AES.r3.t3.t3.s0.clk )
    begin
        case ( \AES.r3.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t3.s4.clk  = \AES.r3.t3.t3.clk ;
    assign \AES.r3.t3.t3.s4.in  = \AES.r3.t3.t3.in ;
    assign \AES.r3.t3.t3.k1  = \AES.r3.t3.t3.s4.out ;
    always @ (  posedge \AES.r3.t3.t3.s4.clk )
    begin
        case ( \AES.r3.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r3.t3.t3.out  = { \AES.r3.t3.t3.k0 , \AES.r3.t3.t3.k0 , ( \AES.r3.t3.t3.k0  ^ \AES.r3.t3.t3.k1  ), \AES.r3.t3.t3.k1  };
    assign \AES.r3.z0  = ( ( ( ( \AES.r3.p00  ^ \AES.r3.p11  ) ^ \AES.r3.p22  ) ^ \AES.r3.p33  ) ^ \AES.r3.k0  );
    assign \AES.r3.z1  = ( ( ( ( \AES.r3.p03  ^ \AES.r3.p10  ) ^ \AES.r3.p21  ) ^ \AES.r3.p32  ) ^ \AES.r3.k1  );
    assign \AES.r3.z2  = ( ( ( ( \AES.r3.p02  ^ \AES.r3.p13  ) ^ \AES.r3.p20  ) ^ \AES.r3.p31  ) ^ \AES.r3.k2  );
    assign \AES.r3.z3  = ( ( ( ( \AES.r3.p01  ^ \AES.r3.p12  ) ^ \AES.r3.p23  ) ^ \AES.r3.p30  ) ^ \AES.r3.k3  );
    always @ (  posedge \AES.r3.clk )
    begin
    end
    assign \AES.r4.clk  = \AES.clk ;
    assign \AES.r4.state_in  = \AES.s3 ;
    assign \AES.r4.key  = \AES.k3b ;
    assign \AES.s4  = \AES.r4.state_out ;
    assign \AES.r4.k0  = \AES.r4.key [127:96];
    assign \AES.r4.k1  = \AES.r4.key [95:64];
    assign \AES.r4.k2  = \AES.r4.key [63:32];
    assign \AES.r4.k3  = \AES.r4.key [31:0];
    assign \AES.r4.s0  = \AES.r4.state_in [127:96];
    assign \AES.r4.s1  = \AES.r4.state_in [95:64];
    assign \AES.r4.s2  = \AES.r4.state_in [63:32];
    assign \AES.r4.s3  = \AES.r4.state_in [31:0];
    assign \AES.r4.t0.clk  = \AES.r4.clk ;
    assign \AES.r4.t0.state  = \AES.r4.s0 ;
    assign \AES.r4.p00  = \AES.r4.t0.p0 ;
    assign \AES.r4.p01  = \AES.r4.t0.p1 ;
    assign \AES.r4.p02  = \AES.r4.t0.p2 ;
    assign \AES.r4.p03  = \AES.r4.t0.p3 ;
    assign \AES.r4.t0.p0  = { \AES.r4.t0.k0 [7:0], \AES.r4.t0.k0 [31:8] };
    assign \AES.r4.t0.p1  = { \AES.r4.t0.k1 [15:0], \AES.r4.t0.k1 [31:16] };
    assign \AES.r4.t0.p2  = { \AES.r4.t0.k2 [23:0], \AES.r4.t0.k2 [31:24] };
    assign \AES.r4.t0.b0  = \AES.r4.t0.state [31:24];
    assign \AES.r4.t0.b1  = \AES.r4.t0.state [23:16];
    assign \AES.r4.t0.b2  = \AES.r4.t0.state [15:8];
    assign \AES.r4.t0.b3  = \AES.r4.t0.state [7:0];
    assign \AES.r4.t0.t0.clk  = \AES.r4.t0.clk ;
    assign \AES.r4.t0.t0.in  = \AES.r4.t0.b0 ;
    assign \AES.r4.t0.k0  = \AES.r4.t0.t0.out ;
    assign \AES.r4.t0.t0.s0.clk  = \AES.r4.t0.t0.clk ;
    assign \AES.r4.t0.t0.s0.in  = \AES.r4.t0.t0.in ;
    assign \AES.r4.t0.t0.k0  = \AES.r4.t0.t0.s0.out ;
    always @ (  posedge \AES.r4.t0.t0.s0.clk )
    begin
        case ( \AES.r4.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t0.s4.clk  = \AES.r4.t0.t0.clk ;
    assign \AES.r4.t0.t0.s4.in  = \AES.r4.t0.t0.in ;
    assign \AES.r4.t0.t0.k1  = \AES.r4.t0.t0.s4.out ;
    always @ (  posedge \AES.r4.t0.t0.s4.clk )
    begin
        case ( \AES.r4.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t0.out  = { \AES.r4.t0.t0.k0 , \AES.r4.t0.t0.k0 , ( \AES.r4.t0.t0.k0  ^ \AES.r4.t0.t0.k1  ), \AES.r4.t0.t0.k1  };
    assign \AES.r4.t0.t1.clk  = \AES.r4.t0.clk ;
    assign \AES.r4.t0.t1.in  = \AES.r4.t0.b1 ;
    assign \AES.r4.t0.k1  = \AES.r4.t0.t1.out ;
    assign \AES.r4.t0.t1.s0.clk  = \AES.r4.t0.t1.clk ;
    assign \AES.r4.t0.t1.s0.in  = \AES.r4.t0.t1.in ;
    assign \AES.r4.t0.t1.k0  = \AES.r4.t0.t1.s0.out ;
    always @ (  posedge \AES.r4.t0.t1.s0.clk )
    begin
        case ( \AES.r4.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t1.s4.clk  = \AES.r4.t0.t1.clk ;
    assign \AES.r4.t0.t1.s4.in  = \AES.r4.t0.t1.in ;
    assign \AES.r4.t0.t1.k1  = \AES.r4.t0.t1.s4.out ;
    always @ (  posedge \AES.r4.t0.t1.s4.clk )
    begin
        case ( \AES.r4.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t1.out  = { \AES.r4.t0.t1.k0 , \AES.r4.t0.t1.k0 , ( \AES.r4.t0.t1.k0  ^ \AES.r4.t0.t1.k1  ), \AES.r4.t0.t1.k1  };
    assign \AES.r4.t0.t2.clk  = \AES.r4.t0.clk ;
    assign \AES.r4.t0.t2.in  = \AES.r4.t0.b2 ;
    assign \AES.r4.t0.k2  = \AES.r4.t0.t2.out ;
    assign \AES.r4.t0.t2.s0.clk  = \AES.r4.t0.t2.clk ;
    assign \AES.r4.t0.t2.s0.in  = \AES.r4.t0.t2.in ;
    assign \AES.r4.t0.t2.k0  = \AES.r4.t0.t2.s0.out ;
    always @ (  posedge \AES.r4.t0.t2.s0.clk )
    begin
        case ( \AES.r4.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t2.s4.clk  = \AES.r4.t0.t2.clk ;
    assign \AES.r4.t0.t2.s4.in  = \AES.r4.t0.t2.in ;
    assign \AES.r4.t0.t2.k1  = \AES.r4.t0.t2.s4.out ;
    always @ (  posedge \AES.r4.t0.t2.s4.clk )
    begin
        case ( \AES.r4.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t2.out  = { \AES.r4.t0.t2.k0 , \AES.r4.t0.t2.k0 , ( \AES.r4.t0.t2.k0  ^ \AES.r4.t0.t2.k1  ), \AES.r4.t0.t2.k1  };
    assign \AES.r4.t0.t3.clk  = \AES.r4.t0.clk ;
    assign \AES.r4.t0.t3.in  = \AES.r4.t0.b3 ;
    assign \AES.r4.t0.p3  = \AES.r4.t0.t3.out ;
    assign \AES.r4.t0.t3.s0.clk  = \AES.r4.t0.t3.clk ;
    assign \AES.r4.t0.t3.s0.in  = \AES.r4.t0.t3.in ;
    assign \AES.r4.t0.t3.k0  = \AES.r4.t0.t3.s0.out ;
    always @ (  posedge \AES.r4.t0.t3.s0.clk )
    begin
        case ( \AES.r4.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t3.s4.clk  = \AES.r4.t0.t3.clk ;
    assign \AES.r4.t0.t3.s4.in  = \AES.r4.t0.t3.in ;
    assign \AES.r4.t0.t3.k1  = \AES.r4.t0.t3.s4.out ;
    always @ (  posedge \AES.r4.t0.t3.s4.clk )
    begin
        case ( \AES.r4.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t0.t3.out  = { \AES.r4.t0.t3.k0 , \AES.r4.t0.t3.k0 , ( \AES.r4.t0.t3.k0  ^ \AES.r4.t0.t3.k1  ), \AES.r4.t0.t3.k1  };
    assign \AES.r4.t1.clk  = \AES.r4.clk ;
    assign \AES.r4.t1.state  = \AES.r4.s1 ;
    assign \AES.r4.p10  = \AES.r4.t1.p0 ;
    assign \AES.r4.p11  = \AES.r4.t1.p1 ;
    assign \AES.r4.p12  = \AES.r4.t1.p2 ;
    assign \AES.r4.p13  = \AES.r4.t1.p3 ;
    assign \AES.r4.t1.p0  = { \AES.r4.t1.k0 [7:0], \AES.r4.t1.k0 [31:8] };
    assign \AES.r4.t1.p1  = { \AES.r4.t1.k1 [15:0], \AES.r4.t1.k1 [31:16] };
    assign \AES.r4.t1.p2  = { \AES.r4.t1.k2 [23:0], \AES.r4.t1.k2 [31:24] };
    assign \AES.r4.t1.b0  = \AES.r4.t1.state [31:24];
    assign \AES.r4.t1.b1  = \AES.r4.t1.state [23:16];
    assign \AES.r4.t1.b2  = \AES.r4.t1.state [15:8];
    assign \AES.r4.t1.b3  = \AES.r4.t1.state [7:0];
    assign \AES.r4.t1.t0.clk  = \AES.r4.t1.clk ;
    assign \AES.r4.t1.t0.in  = \AES.r4.t1.b0 ;
    assign \AES.r4.t1.k0  = \AES.r4.t1.t0.out ;
    assign \AES.r4.t1.t0.s0.clk  = \AES.r4.t1.t0.clk ;
    assign \AES.r4.t1.t0.s0.in  = \AES.r4.t1.t0.in ;
    assign \AES.r4.t1.t0.k0  = \AES.r4.t1.t0.s0.out ;
    always @ (  posedge \AES.r4.t1.t0.s0.clk )
    begin
        case ( \AES.r4.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t0.s4.clk  = \AES.r4.t1.t0.clk ;
    assign \AES.r4.t1.t0.s4.in  = \AES.r4.t1.t0.in ;
    assign \AES.r4.t1.t0.k1  = \AES.r4.t1.t0.s4.out ;
    always @ (  posedge \AES.r4.t1.t0.s4.clk )
    begin
        case ( \AES.r4.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t0.out  = { \AES.r4.t1.t0.k0 , \AES.r4.t1.t0.k0 , ( \AES.r4.t1.t0.k0  ^ \AES.r4.t1.t0.k1  ), \AES.r4.t1.t0.k1  };
    assign \AES.r4.t1.t1.clk  = \AES.r4.t1.clk ;
    assign \AES.r4.t1.t1.in  = \AES.r4.t1.b1 ;
    assign \AES.r4.t1.k1  = \AES.r4.t1.t1.out ;
    assign \AES.r4.t1.t1.s0.clk  = \AES.r4.t1.t1.clk ;
    assign \AES.r4.t1.t1.s0.in  = \AES.r4.t1.t1.in ;
    assign \AES.r4.t1.t1.k0  = \AES.r4.t1.t1.s0.out ;
    always @ (  posedge \AES.r4.t1.t1.s0.clk )
    begin
        case ( \AES.r4.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t1.s4.clk  = \AES.r4.t1.t1.clk ;
    assign \AES.r4.t1.t1.s4.in  = \AES.r4.t1.t1.in ;
    assign \AES.r4.t1.t1.k1  = \AES.r4.t1.t1.s4.out ;
    always @ (  posedge \AES.r4.t1.t1.s4.clk )
    begin
        case ( \AES.r4.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t1.out  = { \AES.r4.t1.t1.k0 , \AES.r4.t1.t1.k0 , ( \AES.r4.t1.t1.k0  ^ \AES.r4.t1.t1.k1  ), \AES.r4.t1.t1.k1  };
    assign \AES.r4.t1.t2.clk  = \AES.r4.t1.clk ;
    assign \AES.r4.t1.t2.in  = \AES.r4.t1.b2 ;
    assign \AES.r4.t1.k2  = \AES.r4.t1.t2.out ;
    assign \AES.r4.t1.t2.s0.clk  = \AES.r4.t1.t2.clk ;
    assign \AES.r4.t1.t2.s0.in  = \AES.r4.t1.t2.in ;
    assign \AES.r4.t1.t2.k0  = \AES.r4.t1.t2.s0.out ;
    always @ (  posedge \AES.r4.t1.t2.s0.clk )
    begin
        case ( \AES.r4.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t2.s4.clk  = \AES.r4.t1.t2.clk ;
    assign \AES.r4.t1.t2.s4.in  = \AES.r4.t1.t2.in ;
    assign \AES.r4.t1.t2.k1  = \AES.r4.t1.t2.s4.out ;
    always @ (  posedge \AES.r4.t1.t2.s4.clk )
    begin
        case ( \AES.r4.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t2.out  = { \AES.r4.t1.t2.k0 , \AES.r4.t1.t2.k0 , ( \AES.r4.t1.t2.k0  ^ \AES.r4.t1.t2.k1  ), \AES.r4.t1.t2.k1  };
    assign \AES.r4.t1.t3.clk  = \AES.r4.t1.clk ;
    assign \AES.r4.t1.t3.in  = \AES.r4.t1.b3 ;
    assign \AES.r4.t1.p3  = \AES.r4.t1.t3.out ;
    assign \AES.r4.t1.t3.s0.clk  = \AES.r4.t1.t3.clk ;
    assign \AES.r4.t1.t3.s0.in  = \AES.r4.t1.t3.in ;
    assign \AES.r4.t1.t3.k0  = \AES.r4.t1.t3.s0.out ;
    always @ (  posedge \AES.r4.t1.t3.s0.clk )
    begin
        case ( \AES.r4.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t3.s4.clk  = \AES.r4.t1.t3.clk ;
    assign \AES.r4.t1.t3.s4.in  = \AES.r4.t1.t3.in ;
    assign \AES.r4.t1.t3.k1  = \AES.r4.t1.t3.s4.out ;
    always @ (  posedge \AES.r4.t1.t3.s4.clk )
    begin
        case ( \AES.r4.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t1.t3.out  = { \AES.r4.t1.t3.k0 , \AES.r4.t1.t3.k0 , ( \AES.r4.t1.t3.k0  ^ \AES.r4.t1.t3.k1  ), \AES.r4.t1.t3.k1  };
    assign \AES.r4.t2.clk  = \AES.r4.clk ;
    assign \AES.r4.t2.state  = \AES.r4.s2 ;
    assign \AES.r4.p20  = \AES.r4.t2.p0 ;
    assign \AES.r4.p21  = \AES.r4.t2.p1 ;
    assign \AES.r4.p22  = \AES.r4.t2.p2 ;
    assign \AES.r4.p23  = \AES.r4.t2.p3 ;
    assign \AES.r4.t2.p0  = { \AES.r4.t2.k0 [7:0], \AES.r4.t2.k0 [31:8] };
    assign \AES.r4.t2.p1  = { \AES.r4.t2.k1 [15:0], \AES.r4.t2.k1 [31:16] };
    assign \AES.r4.t2.p2  = { \AES.r4.t2.k2 [23:0], \AES.r4.t2.k2 [31:24] };
    assign \AES.r4.t2.b0  = \AES.r4.t2.state [31:24];
    assign \AES.r4.t2.b1  = \AES.r4.t2.state [23:16];
    assign \AES.r4.t2.b2  = \AES.r4.t2.state [15:8];
    assign \AES.r4.t2.b3  = \AES.r4.t2.state [7:0];
    assign \AES.r4.t2.t0.clk  = \AES.r4.t2.clk ;
    assign \AES.r4.t2.t0.in  = \AES.r4.t2.b0 ;
    assign \AES.r4.t2.k0  = \AES.r4.t2.t0.out ;
    assign \AES.r4.t2.t0.s0.clk  = \AES.r4.t2.t0.clk ;
    assign \AES.r4.t2.t0.s0.in  = \AES.r4.t2.t0.in ;
    assign \AES.r4.t2.t0.k0  = \AES.r4.t2.t0.s0.out ;
    always @ (  posedge \AES.r4.t2.t0.s0.clk )
    begin
        case ( \AES.r4.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t0.s4.clk  = \AES.r4.t2.t0.clk ;
    assign \AES.r4.t2.t0.s4.in  = \AES.r4.t2.t0.in ;
    assign \AES.r4.t2.t0.k1  = \AES.r4.t2.t0.s4.out ;
    always @ (  posedge \AES.r4.t2.t0.s4.clk )
    begin
        case ( \AES.r4.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t0.out  = { \AES.r4.t2.t0.k0 , \AES.r4.t2.t0.k0 , ( \AES.r4.t2.t0.k0  ^ \AES.r4.t2.t0.k1  ), \AES.r4.t2.t0.k1  };
    assign \AES.r4.t2.t1.clk  = \AES.r4.t2.clk ;
    assign \AES.r4.t2.t1.in  = \AES.r4.t2.b1 ;
    assign \AES.r4.t2.k1  = \AES.r4.t2.t1.out ;
    assign \AES.r4.t2.t1.s0.clk  = \AES.r4.t2.t1.clk ;
    assign \AES.r4.t2.t1.s0.in  = \AES.r4.t2.t1.in ;
    assign \AES.r4.t2.t1.k0  = \AES.r4.t2.t1.s0.out ;
    always @ (  posedge \AES.r4.t2.t1.s0.clk )
    begin
        case ( \AES.r4.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t1.s4.clk  = \AES.r4.t2.t1.clk ;
    assign \AES.r4.t2.t1.s4.in  = \AES.r4.t2.t1.in ;
    assign \AES.r4.t2.t1.k1  = \AES.r4.t2.t1.s4.out ;
    always @ (  posedge \AES.r4.t2.t1.s4.clk )
    begin
        case ( \AES.r4.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t1.out  = { \AES.r4.t2.t1.k0 , \AES.r4.t2.t1.k0 , ( \AES.r4.t2.t1.k0  ^ \AES.r4.t2.t1.k1  ), \AES.r4.t2.t1.k1  };
    assign \AES.r4.t2.t2.clk  = \AES.r4.t2.clk ;
    assign \AES.r4.t2.t2.in  = \AES.r4.t2.b2 ;
    assign \AES.r4.t2.k2  = \AES.r4.t2.t2.out ;
    assign \AES.r4.t2.t2.s0.clk  = \AES.r4.t2.t2.clk ;
    assign \AES.r4.t2.t2.s0.in  = \AES.r4.t2.t2.in ;
    assign \AES.r4.t2.t2.k0  = \AES.r4.t2.t2.s0.out ;
    always @ (  posedge \AES.r4.t2.t2.s0.clk )
    begin
        case ( \AES.r4.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t2.s4.clk  = \AES.r4.t2.t2.clk ;
    assign \AES.r4.t2.t2.s4.in  = \AES.r4.t2.t2.in ;
    assign \AES.r4.t2.t2.k1  = \AES.r4.t2.t2.s4.out ;
    always @ (  posedge \AES.r4.t2.t2.s4.clk )
    begin
        case ( \AES.r4.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t2.out  = { \AES.r4.t2.t2.k0 , \AES.r4.t2.t2.k0 , ( \AES.r4.t2.t2.k0  ^ \AES.r4.t2.t2.k1  ), \AES.r4.t2.t2.k1  };
    assign \AES.r4.t2.t3.clk  = \AES.r4.t2.clk ;
    assign \AES.r4.t2.t3.in  = \AES.r4.t2.b3 ;
    assign \AES.r4.t2.p3  = \AES.r4.t2.t3.out ;
    assign \AES.r4.t2.t3.s0.clk  = \AES.r4.t2.t3.clk ;
    assign \AES.r4.t2.t3.s0.in  = \AES.r4.t2.t3.in ;
    assign \AES.r4.t2.t3.k0  = \AES.r4.t2.t3.s0.out ;
    always @ (  posedge \AES.r4.t2.t3.s0.clk )
    begin
        case ( \AES.r4.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t3.s4.clk  = \AES.r4.t2.t3.clk ;
    assign \AES.r4.t2.t3.s4.in  = \AES.r4.t2.t3.in ;
    assign \AES.r4.t2.t3.k1  = \AES.r4.t2.t3.s4.out ;
    always @ (  posedge \AES.r4.t2.t3.s4.clk )
    begin
        case ( \AES.r4.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t2.t3.out  = { \AES.r4.t2.t3.k0 , \AES.r4.t2.t3.k0 , ( \AES.r4.t2.t3.k0  ^ \AES.r4.t2.t3.k1  ), \AES.r4.t2.t3.k1  };
    assign \AES.r4.t3.clk  = \AES.r4.clk ;
    assign \AES.r4.t3.state  = \AES.r4.s3 ;
    assign \AES.r4.p30  = \AES.r4.t3.p0 ;
    assign \AES.r4.p31  = \AES.r4.t3.p1 ;
    assign \AES.r4.p32  = \AES.r4.t3.p2 ;
    assign \AES.r4.p33  = \AES.r4.t3.p3 ;
    assign \AES.r4.t3.p0  = { \AES.r4.t3.k0 [7:0], \AES.r4.t3.k0 [31:8] };
    assign \AES.r4.t3.p1  = { \AES.r4.t3.k1 [15:0], \AES.r4.t3.k1 [31:16] };
    assign \AES.r4.t3.p2  = { \AES.r4.t3.k2 [23:0], \AES.r4.t3.k2 [31:24] };
    assign \AES.r4.t3.b0  = \AES.r4.t3.state [31:24];
    assign \AES.r4.t3.b1  = \AES.r4.t3.state [23:16];
    assign \AES.r4.t3.b2  = \AES.r4.t3.state [15:8];
    assign \AES.r4.t3.b3  = \AES.r4.t3.state [7:0];
    assign \AES.r4.t3.t0.clk  = \AES.r4.t3.clk ;
    assign \AES.r4.t3.t0.in  = \AES.r4.t3.b0 ;
    assign \AES.r4.t3.k0  = \AES.r4.t3.t0.out ;
    assign \AES.r4.t3.t0.s0.clk  = \AES.r4.t3.t0.clk ;
    assign \AES.r4.t3.t0.s0.in  = \AES.r4.t3.t0.in ;
    assign \AES.r4.t3.t0.k0  = \AES.r4.t3.t0.s0.out ;
    always @ (  posedge \AES.r4.t3.t0.s0.clk )
    begin
        case ( \AES.r4.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t0.s4.clk  = \AES.r4.t3.t0.clk ;
    assign \AES.r4.t3.t0.s4.in  = \AES.r4.t3.t0.in ;
    assign \AES.r4.t3.t0.k1  = \AES.r4.t3.t0.s4.out ;
    always @ (  posedge \AES.r4.t3.t0.s4.clk )
    begin
        case ( \AES.r4.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t0.out  = { \AES.r4.t3.t0.k0 , \AES.r4.t3.t0.k0 , ( \AES.r4.t3.t0.k0  ^ \AES.r4.t3.t0.k1  ), \AES.r4.t3.t0.k1  };
    assign \AES.r4.t3.t1.clk  = \AES.r4.t3.clk ;
    assign \AES.r4.t3.t1.in  = \AES.r4.t3.b1 ;
    assign \AES.r4.t3.k1  = \AES.r4.t3.t1.out ;
    assign \AES.r4.t3.t1.s0.clk  = \AES.r4.t3.t1.clk ;
    assign \AES.r4.t3.t1.s0.in  = \AES.r4.t3.t1.in ;
    assign \AES.r4.t3.t1.k0  = \AES.r4.t3.t1.s0.out ;
    always @ (  posedge \AES.r4.t3.t1.s0.clk )
    begin
        case ( \AES.r4.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t1.s4.clk  = \AES.r4.t3.t1.clk ;
    assign \AES.r4.t3.t1.s4.in  = \AES.r4.t3.t1.in ;
    assign \AES.r4.t3.t1.k1  = \AES.r4.t3.t1.s4.out ;
    always @ (  posedge \AES.r4.t3.t1.s4.clk )
    begin
        case ( \AES.r4.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t1.out  = { \AES.r4.t3.t1.k0 , \AES.r4.t3.t1.k0 , ( \AES.r4.t3.t1.k0  ^ \AES.r4.t3.t1.k1  ), \AES.r4.t3.t1.k1  };
    assign \AES.r4.t3.t2.clk  = \AES.r4.t3.clk ;
    assign \AES.r4.t3.t2.in  = \AES.r4.t3.b2 ;
    assign \AES.r4.t3.k2  = \AES.r4.t3.t2.out ;
    assign \AES.r4.t3.t2.s0.clk  = \AES.r4.t3.t2.clk ;
    assign \AES.r4.t3.t2.s0.in  = \AES.r4.t3.t2.in ;
    assign \AES.r4.t3.t2.k0  = \AES.r4.t3.t2.s0.out ;
    always @ (  posedge \AES.r4.t3.t2.s0.clk )
    begin
        case ( \AES.r4.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t2.s4.clk  = \AES.r4.t3.t2.clk ;
    assign \AES.r4.t3.t2.s4.in  = \AES.r4.t3.t2.in ;
    assign \AES.r4.t3.t2.k1  = \AES.r4.t3.t2.s4.out ;
    always @ (  posedge \AES.r4.t3.t2.s4.clk )
    begin
        case ( \AES.r4.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t2.out  = { \AES.r4.t3.t2.k0 , \AES.r4.t3.t2.k0 , ( \AES.r4.t3.t2.k0  ^ \AES.r4.t3.t2.k1  ), \AES.r4.t3.t2.k1  };
    assign \AES.r4.t3.t3.clk  = \AES.r4.t3.clk ;
    assign \AES.r4.t3.t3.in  = \AES.r4.t3.b3 ;
    assign \AES.r4.t3.p3  = \AES.r4.t3.t3.out ;
    assign \AES.r4.t3.t3.s0.clk  = \AES.r4.t3.t3.clk ;
    assign \AES.r4.t3.t3.s0.in  = \AES.r4.t3.t3.in ;
    assign \AES.r4.t3.t3.k0  = \AES.r4.t3.t3.s0.out ;
    always @ (  posedge \AES.r4.t3.t3.s0.clk )
    begin
        case ( \AES.r4.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t3.s4.clk  = \AES.r4.t3.t3.clk ;
    assign \AES.r4.t3.t3.s4.in  = \AES.r4.t3.t3.in ;
    assign \AES.r4.t3.t3.k1  = \AES.r4.t3.t3.s4.out ;
    always @ (  posedge \AES.r4.t3.t3.s4.clk )
    begin
        case ( \AES.r4.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r4.t3.t3.out  = { \AES.r4.t3.t3.k0 , \AES.r4.t3.t3.k0 , ( \AES.r4.t3.t3.k0  ^ \AES.r4.t3.t3.k1  ), \AES.r4.t3.t3.k1  };
    assign \AES.r4.z0  = ( ( ( ( \AES.r4.p00  ^ \AES.r4.p11  ) ^ \AES.r4.p22  ) ^ \AES.r4.p33  ) ^ \AES.r4.k0  );
    assign \AES.r4.z1  = ( ( ( ( \AES.r4.p03  ^ \AES.r4.p10  ) ^ \AES.r4.p21  ) ^ \AES.r4.p32  ) ^ \AES.r4.k1  );
    assign \AES.r4.z2  = ( ( ( ( \AES.r4.p02  ^ \AES.r4.p13  ) ^ \AES.r4.p20  ) ^ \AES.r4.p31  ) ^ \AES.r4.k2  );
    assign \AES.r4.z3  = ( ( ( ( \AES.r4.p01  ^ \AES.r4.p12  ) ^ \AES.r4.p23  ) ^ \AES.r4.p30  ) ^ \AES.r4.k3  );
    always @ (  posedge \AES.r4.clk )
    begin
    end
    assign \AES.r5.clk  = \AES.clk ;
    assign \AES.r5.state_in  = \AES.s4 ;
    assign \AES.r5.key  = \AES.k4b ;
    assign \AES.s5  = \AES.r5.state_out ;
    assign \AES.r5.k0  = \AES.r5.key [127:96];
    assign \AES.r5.k1  = \AES.r5.key [95:64];
    assign \AES.r5.k2  = \AES.r5.key [63:32];
    assign \AES.r5.k3  = \AES.r5.key [31:0];
    assign \AES.r5.s0  = \AES.r5.state_in [127:96];
    assign \AES.r5.s1  = \AES.r5.state_in [95:64];
    assign \AES.r5.s2  = \AES.r5.state_in [63:32];
    assign \AES.r5.s3  = \AES.r5.state_in [31:0];
    assign \AES.r5.t0.clk  = \AES.r5.clk ;
    assign \AES.r5.t0.state  = \AES.r5.s0 ;
    assign \AES.r5.p00  = \AES.r5.t0.p0 ;
    assign \AES.r5.p01  = \AES.r5.t0.p1 ;
    assign \AES.r5.p02  = \AES.r5.t0.p2 ;
    assign \AES.r5.p03  = \AES.r5.t0.p3 ;
    assign \AES.r5.t0.p0  = { \AES.r5.t0.k0 [7:0], \AES.r5.t0.k0 [31:8] };
    assign \AES.r5.t0.p1  = { \AES.r5.t0.k1 [15:0], \AES.r5.t0.k1 [31:16] };
    assign \AES.r5.t0.p2  = { \AES.r5.t0.k2 [23:0], \AES.r5.t0.k2 [31:24] };
    assign \AES.r5.t0.b0  = \AES.r5.t0.state [31:24];
    assign \AES.r5.t0.b1  = \AES.r5.t0.state [23:16];
    assign \AES.r5.t0.b2  = \AES.r5.t0.state [15:8];
    assign \AES.r5.t0.b3  = \AES.r5.t0.state [7:0];
    assign \AES.r5.t0.t0.clk  = \AES.r5.t0.clk ;
    assign \AES.r5.t0.t0.in  = \AES.r5.t0.b0 ;
    assign \AES.r5.t0.k0  = \AES.r5.t0.t0.out ;
    assign \AES.r5.t0.t0.s0.clk  = \AES.r5.t0.t0.clk ;
    assign \AES.r5.t0.t0.s0.in  = \AES.r5.t0.t0.in ;
    assign \AES.r5.t0.t0.k0  = \AES.r5.t0.t0.s0.out ;
    always @ (  posedge \AES.r5.t0.t0.s0.clk )
    begin
        case ( \AES.r5.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t0.s4.clk  = \AES.r5.t0.t0.clk ;
    assign \AES.r5.t0.t0.s4.in  = \AES.r5.t0.t0.in ;
    assign \AES.r5.t0.t0.k1  = \AES.r5.t0.t0.s4.out ;
    always @ (  posedge \AES.r5.t0.t0.s4.clk )
    begin
        case ( \AES.r5.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t0.out  = { \AES.r5.t0.t0.k0 , \AES.r5.t0.t0.k0 , ( \AES.r5.t0.t0.k0  ^ \AES.r5.t0.t0.k1  ), \AES.r5.t0.t0.k1  };
    assign \AES.r5.t0.t1.clk  = \AES.r5.t0.clk ;
    assign \AES.r5.t0.t1.in  = \AES.r5.t0.b1 ;
    assign \AES.r5.t0.k1  = \AES.r5.t0.t1.out ;
    assign \AES.r5.t0.t1.s0.clk  = \AES.r5.t0.t1.clk ;
    assign \AES.r5.t0.t1.s0.in  = \AES.r5.t0.t1.in ;
    assign \AES.r5.t0.t1.k0  = \AES.r5.t0.t1.s0.out ;
    always @ (  posedge \AES.r5.t0.t1.s0.clk )
    begin
        case ( \AES.r5.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t1.s4.clk  = \AES.r5.t0.t1.clk ;
    assign \AES.r5.t0.t1.s4.in  = \AES.r5.t0.t1.in ;
    assign \AES.r5.t0.t1.k1  = \AES.r5.t0.t1.s4.out ;
    always @ (  posedge \AES.r5.t0.t1.s4.clk )
    begin
        case ( \AES.r5.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t1.out  = { \AES.r5.t0.t1.k0 , \AES.r5.t0.t1.k0 , ( \AES.r5.t0.t1.k0  ^ \AES.r5.t0.t1.k1  ), \AES.r5.t0.t1.k1  };
    assign \AES.r5.t0.t2.clk  = \AES.r5.t0.clk ;
    assign \AES.r5.t0.t2.in  = \AES.r5.t0.b2 ;
    assign \AES.r5.t0.k2  = \AES.r5.t0.t2.out ;
    assign \AES.r5.t0.t2.s0.clk  = \AES.r5.t0.t2.clk ;
    assign \AES.r5.t0.t2.s0.in  = \AES.r5.t0.t2.in ;
    assign \AES.r5.t0.t2.k0  = \AES.r5.t0.t2.s0.out ;
    always @ (  posedge \AES.r5.t0.t2.s0.clk )
    begin
        case ( \AES.r5.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t2.s4.clk  = \AES.r5.t0.t2.clk ;
    assign \AES.r5.t0.t2.s4.in  = \AES.r5.t0.t2.in ;
    assign \AES.r5.t0.t2.k1  = \AES.r5.t0.t2.s4.out ;
    always @ (  posedge \AES.r5.t0.t2.s4.clk )
    begin
        case ( \AES.r5.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t2.out  = { \AES.r5.t0.t2.k0 , \AES.r5.t0.t2.k0 , ( \AES.r5.t0.t2.k0  ^ \AES.r5.t0.t2.k1  ), \AES.r5.t0.t2.k1  };
    assign \AES.r5.t0.t3.clk  = \AES.r5.t0.clk ;
    assign \AES.r5.t0.t3.in  = \AES.r5.t0.b3 ;
    assign \AES.r5.t0.p3  = \AES.r5.t0.t3.out ;
    assign \AES.r5.t0.t3.s0.clk  = \AES.r5.t0.t3.clk ;
    assign \AES.r5.t0.t3.s0.in  = \AES.r5.t0.t3.in ;
    assign \AES.r5.t0.t3.k0  = \AES.r5.t0.t3.s0.out ;
    always @ (  posedge \AES.r5.t0.t3.s0.clk )
    begin
        case ( \AES.r5.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t3.s4.clk  = \AES.r5.t0.t3.clk ;
    assign \AES.r5.t0.t3.s4.in  = \AES.r5.t0.t3.in ;
    assign \AES.r5.t0.t3.k1  = \AES.r5.t0.t3.s4.out ;
    always @ (  posedge \AES.r5.t0.t3.s4.clk )
    begin
        case ( \AES.r5.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t0.t3.out  = { \AES.r5.t0.t3.k0 , \AES.r5.t0.t3.k0 , ( \AES.r5.t0.t3.k0  ^ \AES.r5.t0.t3.k1  ), \AES.r5.t0.t3.k1  };
    assign \AES.r5.t1.clk  = \AES.r5.clk ;
    assign \AES.r5.t1.state  = \AES.r5.s1 ;
    assign \AES.r5.p10  = \AES.r5.t1.p0 ;
    assign \AES.r5.p11  = \AES.r5.t1.p1 ;
    assign \AES.r5.p12  = \AES.r5.t1.p2 ;
    assign \AES.r5.p13  = \AES.r5.t1.p3 ;
    assign \AES.r5.t1.p0  = { \AES.r5.t1.k0 [7:0], \AES.r5.t1.k0 [31:8] };
    assign \AES.r5.t1.p1  = { \AES.r5.t1.k1 [15:0], \AES.r5.t1.k1 [31:16] };
    assign \AES.r5.t1.p2  = { \AES.r5.t1.k2 [23:0], \AES.r5.t1.k2 [31:24] };
    assign \AES.r5.t1.b0  = \AES.r5.t1.state [31:24];
    assign \AES.r5.t1.b1  = \AES.r5.t1.state [23:16];
    assign \AES.r5.t1.b2  = \AES.r5.t1.state [15:8];
    assign \AES.r5.t1.b3  = \AES.r5.t1.state [7:0];
    assign \AES.r5.t1.t0.clk  = \AES.r5.t1.clk ;
    assign \AES.r5.t1.t0.in  = \AES.r5.t1.b0 ;
    assign \AES.r5.t1.k0  = \AES.r5.t1.t0.out ;
    assign \AES.r5.t1.t0.s0.clk  = \AES.r5.t1.t0.clk ;
    assign \AES.r5.t1.t0.s0.in  = \AES.r5.t1.t0.in ;
    assign \AES.r5.t1.t0.k0  = \AES.r5.t1.t0.s0.out ;
    always @ (  posedge \AES.r5.t1.t0.s0.clk )
    begin
        case ( \AES.r5.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t0.s4.clk  = \AES.r5.t1.t0.clk ;
    assign \AES.r5.t1.t0.s4.in  = \AES.r5.t1.t0.in ;
    assign \AES.r5.t1.t0.k1  = \AES.r5.t1.t0.s4.out ;
    always @ (  posedge \AES.r5.t1.t0.s4.clk )
    begin
        case ( \AES.r5.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t0.out  = { \AES.r5.t1.t0.k0 , \AES.r5.t1.t0.k0 , ( \AES.r5.t1.t0.k0  ^ \AES.r5.t1.t0.k1  ), \AES.r5.t1.t0.k1  };
    assign \AES.r5.t1.t1.clk  = \AES.r5.t1.clk ;
    assign \AES.r5.t1.t1.in  = \AES.r5.t1.b1 ;
    assign \AES.r5.t1.k1  = \AES.r5.t1.t1.out ;
    assign \AES.r5.t1.t1.s0.clk  = \AES.r5.t1.t1.clk ;
    assign \AES.r5.t1.t1.s0.in  = \AES.r5.t1.t1.in ;
    assign \AES.r5.t1.t1.k0  = \AES.r5.t1.t1.s0.out ;
    always @ (  posedge \AES.r5.t1.t1.s0.clk )
    begin
        case ( \AES.r5.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t1.s4.clk  = \AES.r5.t1.t1.clk ;
    assign \AES.r5.t1.t1.s4.in  = \AES.r5.t1.t1.in ;
    assign \AES.r5.t1.t1.k1  = \AES.r5.t1.t1.s4.out ;
    always @ (  posedge \AES.r5.t1.t1.s4.clk )
    begin
        case ( \AES.r5.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t1.out  = { \AES.r5.t1.t1.k0 , \AES.r5.t1.t1.k0 , ( \AES.r5.t1.t1.k0  ^ \AES.r5.t1.t1.k1  ), \AES.r5.t1.t1.k1  };
    assign \AES.r5.t1.t2.clk  = \AES.r5.t1.clk ;
    assign \AES.r5.t1.t2.in  = \AES.r5.t1.b2 ;
    assign \AES.r5.t1.k2  = \AES.r5.t1.t2.out ;
    assign \AES.r5.t1.t2.s0.clk  = \AES.r5.t1.t2.clk ;
    assign \AES.r5.t1.t2.s0.in  = \AES.r5.t1.t2.in ;
    assign \AES.r5.t1.t2.k0  = \AES.r5.t1.t2.s0.out ;
    always @ (  posedge \AES.r5.t1.t2.s0.clk )
    begin
        case ( \AES.r5.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t2.s4.clk  = \AES.r5.t1.t2.clk ;
    assign \AES.r5.t1.t2.s4.in  = \AES.r5.t1.t2.in ;
    assign \AES.r5.t1.t2.k1  = \AES.r5.t1.t2.s4.out ;
    always @ (  posedge \AES.r5.t1.t2.s4.clk )
    begin
        case ( \AES.r5.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t2.out  = { \AES.r5.t1.t2.k0 , \AES.r5.t1.t2.k0 , ( \AES.r5.t1.t2.k0  ^ \AES.r5.t1.t2.k1  ), \AES.r5.t1.t2.k1  };
    assign \AES.r5.t1.t3.clk  = \AES.r5.t1.clk ;
    assign \AES.r5.t1.t3.in  = \AES.r5.t1.b3 ;
    assign \AES.r5.t1.p3  = \AES.r5.t1.t3.out ;
    assign \AES.r5.t1.t3.s0.clk  = \AES.r5.t1.t3.clk ;
    assign \AES.r5.t1.t3.s0.in  = \AES.r5.t1.t3.in ;
    assign \AES.r5.t1.t3.k0  = \AES.r5.t1.t3.s0.out ;
    always @ (  posedge \AES.r5.t1.t3.s0.clk )
    begin
        case ( \AES.r5.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t3.s4.clk  = \AES.r5.t1.t3.clk ;
    assign \AES.r5.t1.t3.s4.in  = \AES.r5.t1.t3.in ;
    assign \AES.r5.t1.t3.k1  = \AES.r5.t1.t3.s4.out ;
    always @ (  posedge \AES.r5.t1.t3.s4.clk )
    begin
        case ( \AES.r5.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t1.t3.out  = { \AES.r5.t1.t3.k0 , \AES.r5.t1.t3.k0 , ( \AES.r5.t1.t3.k0  ^ \AES.r5.t1.t3.k1  ), \AES.r5.t1.t3.k1  };
    assign \AES.r5.t2.clk  = \AES.r5.clk ;
    assign \AES.r5.t2.state  = \AES.r5.s2 ;
    assign \AES.r5.p20  = \AES.r5.t2.p0 ;
    assign \AES.r5.p21  = \AES.r5.t2.p1 ;
    assign \AES.r5.p22  = \AES.r5.t2.p2 ;
    assign \AES.r5.p23  = \AES.r5.t2.p3 ;
    assign \AES.r5.t2.p0  = { \AES.r5.t2.k0 [7:0], \AES.r5.t2.k0 [31:8] };
    assign \AES.r5.t2.p1  = { \AES.r5.t2.k1 [15:0], \AES.r5.t2.k1 [31:16] };
    assign \AES.r5.t2.p2  = { \AES.r5.t2.k2 [23:0], \AES.r5.t2.k2 [31:24] };
    assign \AES.r5.t2.b0  = \AES.r5.t2.state [31:24];
    assign \AES.r5.t2.b1  = \AES.r5.t2.state [23:16];
    assign \AES.r5.t2.b2  = \AES.r5.t2.state [15:8];
    assign \AES.r5.t2.b3  = \AES.r5.t2.state [7:0];
    assign \AES.r5.t2.t0.clk  = \AES.r5.t2.clk ;
    assign \AES.r5.t2.t0.in  = \AES.r5.t2.b0 ;
    assign \AES.r5.t2.k0  = \AES.r5.t2.t0.out ;
    assign \AES.r5.t2.t0.s0.clk  = \AES.r5.t2.t0.clk ;
    assign \AES.r5.t2.t0.s0.in  = \AES.r5.t2.t0.in ;
    assign \AES.r5.t2.t0.k0  = \AES.r5.t2.t0.s0.out ;
    always @ (  posedge \AES.r5.t2.t0.s0.clk )
    begin
        case ( \AES.r5.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t0.s4.clk  = \AES.r5.t2.t0.clk ;
    assign \AES.r5.t2.t0.s4.in  = \AES.r5.t2.t0.in ;
    assign \AES.r5.t2.t0.k1  = \AES.r5.t2.t0.s4.out ;
    always @ (  posedge \AES.r5.t2.t0.s4.clk )
    begin
        case ( \AES.r5.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t0.out  = { \AES.r5.t2.t0.k0 , \AES.r5.t2.t0.k0 , ( \AES.r5.t2.t0.k0  ^ \AES.r5.t2.t0.k1  ), \AES.r5.t2.t0.k1  };
    assign \AES.r5.t2.t1.clk  = \AES.r5.t2.clk ;
    assign \AES.r5.t2.t1.in  = \AES.r5.t2.b1 ;
    assign \AES.r5.t2.k1  = \AES.r5.t2.t1.out ;
    assign \AES.r5.t2.t1.s0.clk  = \AES.r5.t2.t1.clk ;
    assign \AES.r5.t2.t1.s0.in  = \AES.r5.t2.t1.in ;
    assign \AES.r5.t2.t1.k0  = \AES.r5.t2.t1.s0.out ;
    always @ (  posedge \AES.r5.t2.t1.s0.clk )
    begin
        case ( \AES.r5.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t1.s4.clk  = \AES.r5.t2.t1.clk ;
    assign \AES.r5.t2.t1.s4.in  = \AES.r5.t2.t1.in ;
    assign \AES.r5.t2.t1.k1  = \AES.r5.t2.t1.s4.out ;
    always @ (  posedge \AES.r5.t2.t1.s4.clk )
    begin
        case ( \AES.r5.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t1.out  = { \AES.r5.t2.t1.k0 , \AES.r5.t2.t1.k0 , ( \AES.r5.t2.t1.k0  ^ \AES.r5.t2.t1.k1  ), \AES.r5.t2.t1.k1  };
    assign \AES.r5.t2.t2.clk  = \AES.r5.t2.clk ;
    assign \AES.r5.t2.t2.in  = \AES.r5.t2.b2 ;
    assign \AES.r5.t2.k2  = \AES.r5.t2.t2.out ;
    assign \AES.r5.t2.t2.s0.clk  = \AES.r5.t2.t2.clk ;
    assign \AES.r5.t2.t2.s0.in  = \AES.r5.t2.t2.in ;
    assign \AES.r5.t2.t2.k0  = \AES.r5.t2.t2.s0.out ;
    always @ (  posedge \AES.r5.t2.t2.s0.clk )
    begin
        case ( \AES.r5.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t2.s4.clk  = \AES.r5.t2.t2.clk ;
    assign \AES.r5.t2.t2.s4.in  = \AES.r5.t2.t2.in ;
    assign \AES.r5.t2.t2.k1  = \AES.r5.t2.t2.s4.out ;
    always @ (  posedge \AES.r5.t2.t2.s4.clk )
    begin
        case ( \AES.r5.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t2.out  = { \AES.r5.t2.t2.k0 , \AES.r5.t2.t2.k0 , ( \AES.r5.t2.t2.k0  ^ \AES.r5.t2.t2.k1  ), \AES.r5.t2.t2.k1  };
    assign \AES.r5.t2.t3.clk  = \AES.r5.t2.clk ;
    assign \AES.r5.t2.t3.in  = \AES.r5.t2.b3 ;
    assign \AES.r5.t2.p3  = \AES.r5.t2.t3.out ;
    assign \AES.r5.t2.t3.s0.clk  = \AES.r5.t2.t3.clk ;
    assign \AES.r5.t2.t3.s0.in  = \AES.r5.t2.t3.in ;
    assign \AES.r5.t2.t3.k0  = \AES.r5.t2.t3.s0.out ;
    always @ (  posedge \AES.r5.t2.t3.s0.clk )
    begin
        case ( \AES.r5.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t3.s4.clk  = \AES.r5.t2.t3.clk ;
    assign \AES.r5.t2.t3.s4.in  = \AES.r5.t2.t3.in ;
    assign \AES.r5.t2.t3.k1  = \AES.r5.t2.t3.s4.out ;
    always @ (  posedge \AES.r5.t2.t3.s4.clk )
    begin
        case ( \AES.r5.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t2.t3.out  = { \AES.r5.t2.t3.k0 , \AES.r5.t2.t3.k0 , ( \AES.r5.t2.t3.k0  ^ \AES.r5.t2.t3.k1  ), \AES.r5.t2.t3.k1  };
    assign \AES.r5.t3.clk  = \AES.r5.clk ;
    assign \AES.r5.t3.state  = \AES.r5.s3 ;
    assign \AES.r5.p30  = \AES.r5.t3.p0 ;
    assign \AES.r5.p31  = \AES.r5.t3.p1 ;
    assign \AES.r5.p32  = \AES.r5.t3.p2 ;
    assign \AES.r5.p33  = \AES.r5.t3.p3 ;
    assign \AES.r5.t3.p0  = { \AES.r5.t3.k0 [7:0], \AES.r5.t3.k0 [31:8] };
    assign \AES.r5.t3.p1  = { \AES.r5.t3.k1 [15:0], \AES.r5.t3.k1 [31:16] };
    assign \AES.r5.t3.p2  = { \AES.r5.t3.k2 [23:0], \AES.r5.t3.k2 [31:24] };
    assign \AES.r5.t3.b0  = \AES.r5.t3.state [31:24];
    assign \AES.r5.t3.b1  = \AES.r5.t3.state [23:16];
    assign \AES.r5.t3.b2  = \AES.r5.t3.state [15:8];
    assign \AES.r5.t3.b3  = \AES.r5.t3.state [7:0];
    assign \AES.r5.t3.t0.clk  = \AES.r5.t3.clk ;
    assign \AES.r5.t3.t0.in  = \AES.r5.t3.b0 ;
    assign \AES.r5.t3.k0  = \AES.r5.t3.t0.out ;
    assign \AES.r5.t3.t0.s0.clk  = \AES.r5.t3.t0.clk ;
    assign \AES.r5.t3.t0.s0.in  = \AES.r5.t3.t0.in ;
    assign \AES.r5.t3.t0.k0  = \AES.r5.t3.t0.s0.out ;
    always @ (  posedge \AES.r5.t3.t0.s0.clk )
    begin
        case ( \AES.r5.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t0.s4.clk  = \AES.r5.t3.t0.clk ;
    assign \AES.r5.t3.t0.s4.in  = \AES.r5.t3.t0.in ;
    assign \AES.r5.t3.t0.k1  = \AES.r5.t3.t0.s4.out ;
    always @ (  posedge \AES.r5.t3.t0.s4.clk )
    begin
        case ( \AES.r5.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t0.out  = { \AES.r5.t3.t0.k0 , \AES.r5.t3.t0.k0 , ( \AES.r5.t3.t0.k0  ^ \AES.r5.t3.t0.k1  ), \AES.r5.t3.t0.k1  };
    assign \AES.r5.t3.t1.clk  = \AES.r5.t3.clk ;
    assign \AES.r5.t3.t1.in  = \AES.r5.t3.b1 ;
    assign \AES.r5.t3.k1  = \AES.r5.t3.t1.out ;
    assign \AES.r5.t3.t1.s0.clk  = \AES.r5.t3.t1.clk ;
    assign \AES.r5.t3.t1.s0.in  = \AES.r5.t3.t1.in ;
    assign \AES.r5.t3.t1.k0  = \AES.r5.t3.t1.s0.out ;
    always @ (  posedge \AES.r5.t3.t1.s0.clk )
    begin
        case ( \AES.r5.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t1.s4.clk  = \AES.r5.t3.t1.clk ;
    assign \AES.r5.t3.t1.s4.in  = \AES.r5.t3.t1.in ;
    assign \AES.r5.t3.t1.k1  = \AES.r5.t3.t1.s4.out ;
    always @ (  posedge \AES.r5.t3.t1.s4.clk )
    begin
        case ( \AES.r5.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t1.out  = { \AES.r5.t3.t1.k0 , \AES.r5.t3.t1.k0 , ( \AES.r5.t3.t1.k0  ^ \AES.r5.t3.t1.k1  ), \AES.r5.t3.t1.k1  };
    assign \AES.r5.t3.t2.clk  = \AES.r5.t3.clk ;
    assign \AES.r5.t3.t2.in  = \AES.r5.t3.b2 ;
    assign \AES.r5.t3.k2  = \AES.r5.t3.t2.out ;
    assign \AES.r5.t3.t2.s0.clk  = \AES.r5.t3.t2.clk ;
    assign \AES.r5.t3.t2.s0.in  = \AES.r5.t3.t2.in ;
    assign \AES.r5.t3.t2.k0  = \AES.r5.t3.t2.s0.out ;
    always @ (  posedge \AES.r5.t3.t2.s0.clk )
    begin
        case ( \AES.r5.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t2.s4.clk  = \AES.r5.t3.t2.clk ;
    assign \AES.r5.t3.t2.s4.in  = \AES.r5.t3.t2.in ;
    assign \AES.r5.t3.t2.k1  = \AES.r5.t3.t2.s4.out ;
    always @ (  posedge \AES.r5.t3.t2.s4.clk )
    begin
        case ( \AES.r5.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t2.out  = { \AES.r5.t3.t2.k0 , \AES.r5.t3.t2.k0 , ( \AES.r5.t3.t2.k0  ^ \AES.r5.t3.t2.k1  ), \AES.r5.t3.t2.k1  };
    assign \AES.r5.t3.t3.clk  = \AES.r5.t3.clk ;
    assign \AES.r5.t3.t3.in  = \AES.r5.t3.b3 ;
    assign \AES.r5.t3.p3  = \AES.r5.t3.t3.out ;
    assign \AES.r5.t3.t3.s0.clk  = \AES.r5.t3.t3.clk ;
    assign \AES.r5.t3.t3.s0.in  = \AES.r5.t3.t3.in ;
    assign \AES.r5.t3.t3.k0  = \AES.r5.t3.t3.s0.out ;
    always @ (  posedge \AES.r5.t3.t3.s0.clk )
    begin
        case ( \AES.r5.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t3.s4.clk  = \AES.r5.t3.t3.clk ;
    assign \AES.r5.t3.t3.s4.in  = \AES.r5.t3.t3.in ;
    assign \AES.r5.t3.t3.k1  = \AES.r5.t3.t3.s4.out ;
    always @ (  posedge \AES.r5.t3.t3.s4.clk )
    begin
        case ( \AES.r5.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r5.t3.t3.out  = { \AES.r5.t3.t3.k0 , \AES.r5.t3.t3.k0 , ( \AES.r5.t3.t3.k0  ^ \AES.r5.t3.t3.k1  ), \AES.r5.t3.t3.k1  };
    assign \AES.r5.z0  = ( ( ( ( \AES.r5.p00  ^ \AES.r5.p11  ) ^ \AES.r5.p22  ) ^ \AES.r5.p33  ) ^ \AES.r5.k0  );
    assign \AES.r5.z1  = ( ( ( ( \AES.r5.p03  ^ \AES.r5.p10  ) ^ \AES.r5.p21  ) ^ \AES.r5.p32  ) ^ \AES.r5.k1  );
    assign \AES.r5.z2  = ( ( ( ( \AES.r5.p02  ^ \AES.r5.p13  ) ^ \AES.r5.p20  ) ^ \AES.r5.p31  ) ^ \AES.r5.k2  );
    assign \AES.r5.z3  = ( ( ( ( \AES.r5.p01  ^ \AES.r5.p12  ) ^ \AES.r5.p23  ) ^ \AES.r5.p30  ) ^ \AES.r5.k3  );
    always @ (  posedge \AES.r5.clk )
    begin
    end
    assign \AES.r6.clk  = \AES.clk ;
    assign \AES.r6.state_in  = \AES.s5 ;
    assign \AES.r6.key  = \AES.k5b ;
    assign \AES.s6  = \AES.r6.state_out ;
    assign \AES.r6.k0  = \AES.r6.key [127:96];
    assign \AES.r6.k1  = \AES.r6.key [95:64];
    assign \AES.r6.k2  = \AES.r6.key [63:32];
    assign \AES.r6.k3  = \AES.r6.key [31:0];
    assign \AES.r6.s0  = \AES.r6.state_in [127:96];
    assign \AES.r6.s1  = \AES.r6.state_in [95:64];
    assign \AES.r6.s2  = \AES.r6.state_in [63:32];
    assign \AES.r6.s3  = \AES.r6.state_in [31:0];
    assign \AES.r6.t0.clk  = \AES.r6.clk ;
    assign \AES.r6.t0.state  = \AES.r6.s0 ;
    assign \AES.r6.p00  = \AES.r6.t0.p0 ;
    assign \AES.r6.p01  = \AES.r6.t0.p1 ;
    assign \AES.r6.p02  = \AES.r6.t0.p2 ;
    assign \AES.r6.p03  = \AES.r6.t0.p3 ;
    assign \AES.r6.t0.p0  = { \AES.r6.t0.k0 [7:0], \AES.r6.t0.k0 [31:8] };
    assign \AES.r6.t0.p1  = { \AES.r6.t0.k1 [15:0], \AES.r6.t0.k1 [31:16] };
    assign \AES.r6.t0.p2  = { \AES.r6.t0.k2 [23:0], \AES.r6.t0.k2 [31:24] };
    assign \AES.r6.t0.b0  = \AES.r6.t0.state [31:24];
    assign \AES.r6.t0.b1  = \AES.r6.t0.state [23:16];
    assign \AES.r6.t0.b2  = \AES.r6.t0.state [15:8];
    assign \AES.r6.t0.b3  = \AES.r6.t0.state [7:0];
    assign \AES.r6.t0.t0.clk  = \AES.r6.t0.clk ;
    assign \AES.r6.t0.t0.in  = \AES.r6.t0.b0 ;
    assign \AES.r6.t0.k0  = \AES.r6.t0.t0.out ;
    assign \AES.r6.t0.t0.s0.clk  = \AES.r6.t0.t0.clk ;
    assign \AES.r6.t0.t0.s0.in  = \AES.r6.t0.t0.in ;
    assign \AES.r6.t0.t0.k0  = \AES.r6.t0.t0.s0.out ;
    always @ (  posedge \AES.r6.t0.t0.s0.clk )
    begin
        case ( \AES.r6.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t0.s4.clk  = \AES.r6.t0.t0.clk ;
    assign \AES.r6.t0.t0.s4.in  = \AES.r6.t0.t0.in ;
    assign \AES.r6.t0.t0.k1  = \AES.r6.t0.t0.s4.out ;
    always @ (  posedge \AES.r6.t0.t0.s4.clk )
    begin
        case ( \AES.r6.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t0.out  = { \AES.r6.t0.t0.k0 , \AES.r6.t0.t0.k0 , ( \AES.r6.t0.t0.k0  ^ \AES.r6.t0.t0.k1  ), \AES.r6.t0.t0.k1  };
    assign \AES.r6.t0.t1.clk  = \AES.r6.t0.clk ;
    assign \AES.r6.t0.t1.in  = \AES.r6.t0.b1 ;
    assign \AES.r6.t0.k1  = \AES.r6.t0.t1.out ;
    assign \AES.r6.t0.t1.s0.clk  = \AES.r6.t0.t1.clk ;
    assign \AES.r6.t0.t1.s0.in  = \AES.r6.t0.t1.in ;
    assign \AES.r6.t0.t1.k0  = \AES.r6.t0.t1.s0.out ;
    always @ (  posedge \AES.r6.t0.t1.s0.clk )
    begin
        case ( \AES.r6.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t1.s4.clk  = \AES.r6.t0.t1.clk ;
    assign \AES.r6.t0.t1.s4.in  = \AES.r6.t0.t1.in ;
    assign \AES.r6.t0.t1.k1  = \AES.r6.t0.t1.s4.out ;
    always @ (  posedge \AES.r6.t0.t1.s4.clk )
    begin
        case ( \AES.r6.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t1.out  = { \AES.r6.t0.t1.k0 , \AES.r6.t0.t1.k0 , ( \AES.r6.t0.t1.k0  ^ \AES.r6.t0.t1.k1  ), \AES.r6.t0.t1.k1  };
    assign \AES.r6.t0.t2.clk  = \AES.r6.t0.clk ;
    assign \AES.r6.t0.t2.in  = \AES.r6.t0.b2 ;
    assign \AES.r6.t0.k2  = \AES.r6.t0.t2.out ;
    assign \AES.r6.t0.t2.s0.clk  = \AES.r6.t0.t2.clk ;
    assign \AES.r6.t0.t2.s0.in  = \AES.r6.t0.t2.in ;
    assign \AES.r6.t0.t2.k0  = \AES.r6.t0.t2.s0.out ;
    always @ (  posedge \AES.r6.t0.t2.s0.clk )
    begin
        case ( \AES.r6.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t2.s4.clk  = \AES.r6.t0.t2.clk ;
    assign \AES.r6.t0.t2.s4.in  = \AES.r6.t0.t2.in ;
    assign \AES.r6.t0.t2.k1  = \AES.r6.t0.t2.s4.out ;
    always @ (  posedge \AES.r6.t0.t2.s4.clk )
    begin
        case ( \AES.r6.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t2.out  = { \AES.r6.t0.t2.k0 , \AES.r6.t0.t2.k0 , ( \AES.r6.t0.t2.k0  ^ \AES.r6.t0.t2.k1  ), \AES.r6.t0.t2.k1  };
    assign \AES.r6.t0.t3.clk  = \AES.r6.t0.clk ;
    assign \AES.r6.t0.t3.in  = \AES.r6.t0.b3 ;
    assign \AES.r6.t0.p3  = \AES.r6.t0.t3.out ;
    assign \AES.r6.t0.t3.s0.clk  = \AES.r6.t0.t3.clk ;
    assign \AES.r6.t0.t3.s0.in  = \AES.r6.t0.t3.in ;
    assign \AES.r6.t0.t3.k0  = \AES.r6.t0.t3.s0.out ;
    always @ (  posedge \AES.r6.t0.t3.s0.clk )
    begin
        case ( \AES.r6.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t3.s4.clk  = \AES.r6.t0.t3.clk ;
    assign \AES.r6.t0.t3.s4.in  = \AES.r6.t0.t3.in ;
    assign \AES.r6.t0.t3.k1  = \AES.r6.t0.t3.s4.out ;
    always @ (  posedge \AES.r6.t0.t3.s4.clk )
    begin
        case ( \AES.r6.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t0.t3.out  = { \AES.r6.t0.t3.k0 , \AES.r6.t0.t3.k0 , ( \AES.r6.t0.t3.k0  ^ \AES.r6.t0.t3.k1  ), \AES.r6.t0.t3.k1  };
    assign \AES.r6.t1.clk  = \AES.r6.clk ;
    assign \AES.r6.t1.state  = \AES.r6.s1 ;
    assign \AES.r6.p10  = \AES.r6.t1.p0 ;
    assign \AES.r6.p11  = \AES.r6.t1.p1 ;
    assign \AES.r6.p12  = \AES.r6.t1.p2 ;
    assign \AES.r6.p13  = \AES.r6.t1.p3 ;
    assign \AES.r6.t1.p0  = { \AES.r6.t1.k0 [7:0], \AES.r6.t1.k0 [31:8] };
    assign \AES.r6.t1.p1  = { \AES.r6.t1.k1 [15:0], \AES.r6.t1.k1 [31:16] };
    assign \AES.r6.t1.p2  = { \AES.r6.t1.k2 [23:0], \AES.r6.t1.k2 [31:24] };
    assign \AES.r6.t1.b0  = \AES.r6.t1.state [31:24];
    assign \AES.r6.t1.b1  = \AES.r6.t1.state [23:16];
    assign \AES.r6.t1.b2  = \AES.r6.t1.state [15:8];
    assign \AES.r6.t1.b3  = \AES.r6.t1.state [7:0];
    assign \AES.r6.t1.t0.clk  = \AES.r6.t1.clk ;
    assign \AES.r6.t1.t0.in  = \AES.r6.t1.b0 ;
    assign \AES.r6.t1.k0  = \AES.r6.t1.t0.out ;
    assign \AES.r6.t1.t0.s0.clk  = \AES.r6.t1.t0.clk ;
    assign \AES.r6.t1.t0.s0.in  = \AES.r6.t1.t0.in ;
    assign \AES.r6.t1.t0.k0  = \AES.r6.t1.t0.s0.out ;
    always @ (  posedge \AES.r6.t1.t0.s0.clk )
    begin
        case ( \AES.r6.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t0.s4.clk  = \AES.r6.t1.t0.clk ;
    assign \AES.r6.t1.t0.s4.in  = \AES.r6.t1.t0.in ;
    assign \AES.r6.t1.t0.k1  = \AES.r6.t1.t0.s4.out ;
    always @ (  posedge \AES.r6.t1.t0.s4.clk )
    begin
        case ( \AES.r6.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t0.out  = { \AES.r6.t1.t0.k0 , \AES.r6.t1.t0.k0 , ( \AES.r6.t1.t0.k0  ^ \AES.r6.t1.t0.k1  ), \AES.r6.t1.t0.k1  };
    assign \AES.r6.t1.t1.clk  = \AES.r6.t1.clk ;
    assign \AES.r6.t1.t1.in  = \AES.r6.t1.b1 ;
    assign \AES.r6.t1.k1  = \AES.r6.t1.t1.out ;
    assign \AES.r6.t1.t1.s0.clk  = \AES.r6.t1.t1.clk ;
    assign \AES.r6.t1.t1.s0.in  = \AES.r6.t1.t1.in ;
    assign \AES.r6.t1.t1.k0  = \AES.r6.t1.t1.s0.out ;
    always @ (  posedge \AES.r6.t1.t1.s0.clk )
    begin
        case ( \AES.r6.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t1.s4.clk  = \AES.r6.t1.t1.clk ;
    assign \AES.r6.t1.t1.s4.in  = \AES.r6.t1.t1.in ;
    assign \AES.r6.t1.t1.k1  = \AES.r6.t1.t1.s4.out ;
    always @ (  posedge \AES.r6.t1.t1.s4.clk )
    begin
        case ( \AES.r6.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t1.out  = { \AES.r6.t1.t1.k0 , \AES.r6.t1.t1.k0 , ( \AES.r6.t1.t1.k0  ^ \AES.r6.t1.t1.k1  ), \AES.r6.t1.t1.k1  };
    assign \AES.r6.t1.t2.clk  = \AES.r6.t1.clk ;
    assign \AES.r6.t1.t2.in  = \AES.r6.t1.b2 ;
    assign \AES.r6.t1.k2  = \AES.r6.t1.t2.out ;
    assign \AES.r6.t1.t2.s0.clk  = \AES.r6.t1.t2.clk ;
    assign \AES.r6.t1.t2.s0.in  = \AES.r6.t1.t2.in ;
    assign \AES.r6.t1.t2.k0  = \AES.r6.t1.t2.s0.out ;
    always @ (  posedge \AES.r6.t1.t2.s0.clk )
    begin
        case ( \AES.r6.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t2.s4.clk  = \AES.r6.t1.t2.clk ;
    assign \AES.r6.t1.t2.s4.in  = \AES.r6.t1.t2.in ;
    assign \AES.r6.t1.t2.k1  = \AES.r6.t1.t2.s4.out ;
    always @ (  posedge \AES.r6.t1.t2.s4.clk )
    begin
        case ( \AES.r6.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t2.out  = { \AES.r6.t1.t2.k0 , \AES.r6.t1.t2.k0 , ( \AES.r6.t1.t2.k0  ^ \AES.r6.t1.t2.k1  ), \AES.r6.t1.t2.k1  };
    assign \AES.r6.t1.t3.clk  = \AES.r6.t1.clk ;
    assign \AES.r6.t1.t3.in  = \AES.r6.t1.b3 ;
    assign \AES.r6.t1.p3  = \AES.r6.t1.t3.out ;
    assign \AES.r6.t1.t3.s0.clk  = \AES.r6.t1.t3.clk ;
    assign \AES.r6.t1.t3.s0.in  = \AES.r6.t1.t3.in ;
    assign \AES.r6.t1.t3.k0  = \AES.r6.t1.t3.s0.out ;
    always @ (  posedge \AES.r6.t1.t3.s0.clk )
    begin
        case ( \AES.r6.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t3.s4.clk  = \AES.r6.t1.t3.clk ;
    assign \AES.r6.t1.t3.s4.in  = \AES.r6.t1.t3.in ;
    assign \AES.r6.t1.t3.k1  = \AES.r6.t1.t3.s4.out ;
    always @ (  posedge \AES.r6.t1.t3.s4.clk )
    begin
        case ( \AES.r6.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t1.t3.out  = { \AES.r6.t1.t3.k0 , \AES.r6.t1.t3.k0 , ( \AES.r6.t1.t3.k0  ^ \AES.r6.t1.t3.k1  ), \AES.r6.t1.t3.k1  };
    assign \AES.r6.t2.clk  = \AES.r6.clk ;
    assign \AES.r6.t2.state  = \AES.r6.s2 ;
    assign \AES.r6.p20  = \AES.r6.t2.p0 ;
    assign \AES.r6.p21  = \AES.r6.t2.p1 ;
    assign \AES.r6.p22  = \AES.r6.t2.p2 ;
    assign \AES.r6.p23  = \AES.r6.t2.p3 ;
    assign \AES.r6.t2.p0  = { \AES.r6.t2.k0 [7:0], \AES.r6.t2.k0 [31:8] };
    assign \AES.r6.t2.p1  = { \AES.r6.t2.k1 [15:0], \AES.r6.t2.k1 [31:16] };
    assign \AES.r6.t2.p2  = { \AES.r6.t2.k2 [23:0], \AES.r6.t2.k2 [31:24] };
    assign \AES.r6.t2.b0  = \AES.r6.t2.state [31:24];
    assign \AES.r6.t2.b1  = \AES.r6.t2.state [23:16];
    assign \AES.r6.t2.b2  = \AES.r6.t2.state [15:8];
    assign \AES.r6.t2.b3  = \AES.r6.t2.state [7:0];
    assign \AES.r6.t2.t0.clk  = \AES.r6.t2.clk ;
    assign \AES.r6.t2.t0.in  = \AES.r6.t2.b0 ;
    assign \AES.r6.t2.k0  = \AES.r6.t2.t0.out ;
    assign \AES.r6.t2.t0.s0.clk  = \AES.r6.t2.t0.clk ;
    assign \AES.r6.t2.t0.s0.in  = \AES.r6.t2.t0.in ;
    assign \AES.r6.t2.t0.k0  = \AES.r6.t2.t0.s0.out ;
    always @ (  posedge \AES.r6.t2.t0.s0.clk )
    begin
        case ( \AES.r6.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t0.s4.clk  = \AES.r6.t2.t0.clk ;
    assign \AES.r6.t2.t0.s4.in  = \AES.r6.t2.t0.in ;
    assign \AES.r6.t2.t0.k1  = \AES.r6.t2.t0.s4.out ;
    always @ (  posedge \AES.r6.t2.t0.s4.clk )
    begin
        case ( \AES.r6.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t0.out  = { \AES.r6.t2.t0.k0 , \AES.r6.t2.t0.k0 , ( \AES.r6.t2.t0.k0  ^ \AES.r6.t2.t0.k1  ), \AES.r6.t2.t0.k1  };
    assign \AES.r6.t2.t1.clk  = \AES.r6.t2.clk ;
    assign \AES.r6.t2.t1.in  = \AES.r6.t2.b1 ;
    assign \AES.r6.t2.k1  = \AES.r6.t2.t1.out ;
    assign \AES.r6.t2.t1.s0.clk  = \AES.r6.t2.t1.clk ;
    assign \AES.r6.t2.t1.s0.in  = \AES.r6.t2.t1.in ;
    assign \AES.r6.t2.t1.k0  = \AES.r6.t2.t1.s0.out ;
    always @ (  posedge \AES.r6.t2.t1.s0.clk )
    begin
        case ( \AES.r6.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t1.s4.clk  = \AES.r6.t2.t1.clk ;
    assign \AES.r6.t2.t1.s4.in  = \AES.r6.t2.t1.in ;
    assign \AES.r6.t2.t1.k1  = \AES.r6.t2.t1.s4.out ;
    always @ (  posedge \AES.r6.t2.t1.s4.clk )
    begin
        case ( \AES.r6.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t1.out  = { \AES.r6.t2.t1.k0 , \AES.r6.t2.t1.k0 , ( \AES.r6.t2.t1.k0  ^ \AES.r6.t2.t1.k1  ), \AES.r6.t2.t1.k1  };
    assign \AES.r6.t2.t2.clk  = \AES.r6.t2.clk ;
    assign \AES.r6.t2.t2.in  = \AES.r6.t2.b2 ;
    assign \AES.r6.t2.k2  = \AES.r6.t2.t2.out ;
    assign \AES.r6.t2.t2.s0.clk  = \AES.r6.t2.t2.clk ;
    assign \AES.r6.t2.t2.s0.in  = \AES.r6.t2.t2.in ;
    assign \AES.r6.t2.t2.k0  = \AES.r6.t2.t2.s0.out ;
    always @ (  posedge \AES.r6.t2.t2.s0.clk )
    begin
        case ( \AES.r6.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t2.s4.clk  = \AES.r6.t2.t2.clk ;
    assign \AES.r6.t2.t2.s4.in  = \AES.r6.t2.t2.in ;
    assign \AES.r6.t2.t2.k1  = \AES.r6.t2.t2.s4.out ;
    always @ (  posedge \AES.r6.t2.t2.s4.clk )
    begin
        case ( \AES.r6.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t2.out  = { \AES.r6.t2.t2.k0 , \AES.r6.t2.t2.k0 , ( \AES.r6.t2.t2.k0  ^ \AES.r6.t2.t2.k1  ), \AES.r6.t2.t2.k1  };
    assign \AES.r6.t2.t3.clk  = \AES.r6.t2.clk ;
    assign \AES.r6.t2.t3.in  = \AES.r6.t2.b3 ;
    assign \AES.r6.t2.p3  = \AES.r6.t2.t3.out ;
    assign \AES.r6.t2.t3.s0.clk  = \AES.r6.t2.t3.clk ;
    assign \AES.r6.t2.t3.s0.in  = \AES.r6.t2.t3.in ;
    assign \AES.r6.t2.t3.k0  = \AES.r6.t2.t3.s0.out ;
    always @ (  posedge \AES.r6.t2.t3.s0.clk )
    begin
        case ( \AES.r6.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t3.s4.clk  = \AES.r6.t2.t3.clk ;
    assign \AES.r6.t2.t3.s4.in  = \AES.r6.t2.t3.in ;
    assign \AES.r6.t2.t3.k1  = \AES.r6.t2.t3.s4.out ;
    always @ (  posedge \AES.r6.t2.t3.s4.clk )
    begin
        case ( \AES.r6.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t2.t3.out  = { \AES.r6.t2.t3.k0 , \AES.r6.t2.t3.k0 , ( \AES.r6.t2.t3.k0  ^ \AES.r6.t2.t3.k1  ), \AES.r6.t2.t3.k1  };
    assign \AES.r6.t3.clk  = \AES.r6.clk ;
    assign \AES.r6.t3.state  = \AES.r6.s3 ;
    assign \AES.r6.p30  = \AES.r6.t3.p0 ;
    assign \AES.r6.p31  = \AES.r6.t3.p1 ;
    assign \AES.r6.p32  = \AES.r6.t3.p2 ;
    assign \AES.r6.p33  = \AES.r6.t3.p3 ;
    assign \AES.r6.t3.p0  = { \AES.r6.t3.k0 [7:0], \AES.r6.t3.k0 [31:8] };
    assign \AES.r6.t3.p1  = { \AES.r6.t3.k1 [15:0], \AES.r6.t3.k1 [31:16] };
    assign \AES.r6.t3.p2  = { \AES.r6.t3.k2 [23:0], \AES.r6.t3.k2 [31:24] };
    assign \AES.r6.t3.b0  = \AES.r6.t3.state [31:24];
    assign \AES.r6.t3.b1  = \AES.r6.t3.state [23:16];
    assign \AES.r6.t3.b2  = \AES.r6.t3.state [15:8];
    assign \AES.r6.t3.b3  = \AES.r6.t3.state [7:0];
    assign \AES.r6.t3.t0.clk  = \AES.r6.t3.clk ;
    assign \AES.r6.t3.t0.in  = \AES.r6.t3.b0 ;
    assign \AES.r6.t3.k0  = \AES.r6.t3.t0.out ;
    assign \AES.r6.t3.t0.s0.clk  = \AES.r6.t3.t0.clk ;
    assign \AES.r6.t3.t0.s0.in  = \AES.r6.t3.t0.in ;
    assign \AES.r6.t3.t0.k0  = \AES.r6.t3.t0.s0.out ;
    always @ (  posedge \AES.r6.t3.t0.s0.clk )
    begin
        case ( \AES.r6.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t0.s4.clk  = \AES.r6.t3.t0.clk ;
    assign \AES.r6.t3.t0.s4.in  = \AES.r6.t3.t0.in ;
    assign \AES.r6.t3.t0.k1  = \AES.r6.t3.t0.s4.out ;
    always @ (  posedge \AES.r6.t3.t0.s4.clk )
    begin
        case ( \AES.r6.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t0.out  = { \AES.r6.t3.t0.k0 , \AES.r6.t3.t0.k0 , ( \AES.r6.t3.t0.k0  ^ \AES.r6.t3.t0.k1  ), \AES.r6.t3.t0.k1  };
    assign \AES.r6.t3.t1.clk  = \AES.r6.t3.clk ;
    assign \AES.r6.t3.t1.in  = \AES.r6.t3.b1 ;
    assign \AES.r6.t3.k1  = \AES.r6.t3.t1.out ;
    assign \AES.r6.t3.t1.s0.clk  = \AES.r6.t3.t1.clk ;
    assign \AES.r6.t3.t1.s0.in  = \AES.r6.t3.t1.in ;
    assign \AES.r6.t3.t1.k0  = \AES.r6.t3.t1.s0.out ;
    always @ (  posedge \AES.r6.t3.t1.s0.clk )
    begin
        case ( \AES.r6.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t1.s4.clk  = \AES.r6.t3.t1.clk ;
    assign \AES.r6.t3.t1.s4.in  = \AES.r6.t3.t1.in ;
    assign \AES.r6.t3.t1.k1  = \AES.r6.t3.t1.s4.out ;
    always @ (  posedge \AES.r6.t3.t1.s4.clk )
    begin
        case ( \AES.r6.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t1.out  = { \AES.r6.t3.t1.k0 , \AES.r6.t3.t1.k0 , ( \AES.r6.t3.t1.k0  ^ \AES.r6.t3.t1.k1  ), \AES.r6.t3.t1.k1  };
    assign \AES.r6.t3.t2.clk  = \AES.r6.t3.clk ;
    assign \AES.r6.t3.t2.in  = \AES.r6.t3.b2 ;
    assign \AES.r6.t3.k2  = \AES.r6.t3.t2.out ;
    assign \AES.r6.t3.t2.s0.clk  = \AES.r6.t3.t2.clk ;
    assign \AES.r6.t3.t2.s0.in  = \AES.r6.t3.t2.in ;
    assign \AES.r6.t3.t2.k0  = \AES.r6.t3.t2.s0.out ;
    always @ (  posedge \AES.r6.t3.t2.s0.clk )
    begin
        case ( \AES.r6.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t2.s4.clk  = \AES.r6.t3.t2.clk ;
    assign \AES.r6.t3.t2.s4.in  = \AES.r6.t3.t2.in ;
    assign \AES.r6.t3.t2.k1  = \AES.r6.t3.t2.s4.out ;
    always @ (  posedge \AES.r6.t3.t2.s4.clk )
    begin
        case ( \AES.r6.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t2.out  = { \AES.r6.t3.t2.k0 , \AES.r6.t3.t2.k0 , ( \AES.r6.t3.t2.k0  ^ \AES.r6.t3.t2.k1  ), \AES.r6.t3.t2.k1  };
    assign \AES.r6.t3.t3.clk  = \AES.r6.t3.clk ;
    assign \AES.r6.t3.t3.in  = \AES.r6.t3.b3 ;
    assign \AES.r6.t3.p3  = \AES.r6.t3.t3.out ;
    assign \AES.r6.t3.t3.s0.clk  = \AES.r6.t3.t3.clk ;
    assign \AES.r6.t3.t3.s0.in  = \AES.r6.t3.t3.in ;
    assign \AES.r6.t3.t3.k0  = \AES.r6.t3.t3.s0.out ;
    always @ (  posedge \AES.r6.t3.t3.s0.clk )
    begin
        case ( \AES.r6.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t3.s4.clk  = \AES.r6.t3.t3.clk ;
    assign \AES.r6.t3.t3.s4.in  = \AES.r6.t3.t3.in ;
    assign \AES.r6.t3.t3.k1  = \AES.r6.t3.t3.s4.out ;
    always @ (  posedge \AES.r6.t3.t3.s4.clk )
    begin
        case ( \AES.r6.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r6.t3.t3.out  = { \AES.r6.t3.t3.k0 , \AES.r6.t3.t3.k0 , ( \AES.r6.t3.t3.k0  ^ \AES.r6.t3.t3.k1  ), \AES.r6.t3.t3.k1  };
    assign \AES.r6.z0  = ( ( ( ( \AES.r6.p00  ^ \AES.r6.p11  ) ^ \AES.r6.p22  ) ^ \AES.r6.p33  ) ^ \AES.r6.k0  );
    assign \AES.r6.z1  = ( ( ( ( \AES.r6.p03  ^ \AES.r6.p10  ) ^ \AES.r6.p21  ) ^ \AES.r6.p32  ) ^ \AES.r6.k1  );
    assign \AES.r6.z2  = ( ( ( ( \AES.r6.p02  ^ \AES.r6.p13  ) ^ \AES.r6.p20  ) ^ \AES.r6.p31  ) ^ \AES.r6.k2  );
    assign \AES.r6.z3  = ( ( ( ( \AES.r6.p01  ^ \AES.r6.p12  ) ^ \AES.r6.p23  ) ^ \AES.r6.p30  ) ^ \AES.r6.k3  );
    always @ (  posedge \AES.r6.clk )
    begin
    end
    assign \AES.r7.clk  = \AES.clk ;
    assign \AES.r7.state_in  = \AES.s6 ;
    assign \AES.r7.key  = \AES.k6b ;
    assign \AES.s7  = \AES.r7.state_out ;
    assign \AES.r7.k0  = \AES.r7.key [127:96];
    assign \AES.r7.k1  = \AES.r7.key [95:64];
    assign \AES.r7.k2  = \AES.r7.key [63:32];
    assign \AES.r7.k3  = \AES.r7.key [31:0];
    assign \AES.r7.s0  = \AES.r7.state_in [127:96];
    assign \AES.r7.s1  = \AES.r7.state_in [95:64];
    assign \AES.r7.s2  = \AES.r7.state_in [63:32];
    assign \AES.r7.s3  = \AES.r7.state_in [31:0];
    assign \AES.r7.t0.clk  = \AES.r7.clk ;
    assign \AES.r7.t0.state  = \AES.r7.s0 ;
    assign \AES.r7.p00  = \AES.r7.t0.p0 ;
    assign \AES.r7.p01  = \AES.r7.t0.p1 ;
    assign \AES.r7.p02  = \AES.r7.t0.p2 ;
    assign \AES.r7.p03  = \AES.r7.t0.p3 ;
    assign \AES.r7.t0.p0  = { \AES.r7.t0.k0 [7:0], \AES.r7.t0.k0 [31:8] };
    assign \AES.r7.t0.p1  = { \AES.r7.t0.k1 [15:0], \AES.r7.t0.k1 [31:16] };
    assign \AES.r7.t0.p2  = { \AES.r7.t0.k2 [23:0], \AES.r7.t0.k2 [31:24] };
    assign \AES.r7.t0.b0  = \AES.r7.t0.state [31:24];
    assign \AES.r7.t0.b1  = \AES.r7.t0.state [23:16];
    assign \AES.r7.t0.b2  = \AES.r7.t0.state [15:8];
    assign \AES.r7.t0.b3  = \AES.r7.t0.state [7:0];
    assign \AES.r7.t0.t0.clk  = \AES.r7.t0.clk ;
    assign \AES.r7.t0.t0.in  = \AES.r7.t0.b0 ;
    assign \AES.r7.t0.k0  = \AES.r7.t0.t0.out ;
    assign \AES.r7.t0.t0.s0.clk  = \AES.r7.t0.t0.clk ;
    assign \AES.r7.t0.t0.s0.in  = \AES.r7.t0.t0.in ;
    assign \AES.r7.t0.t0.k0  = \AES.r7.t0.t0.s0.out ;
    always @ (  posedge \AES.r7.t0.t0.s0.clk )
    begin
        case ( \AES.r7.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t0.s4.clk  = \AES.r7.t0.t0.clk ;
    assign \AES.r7.t0.t0.s4.in  = \AES.r7.t0.t0.in ;
    assign \AES.r7.t0.t0.k1  = \AES.r7.t0.t0.s4.out ;
    always @ (  posedge \AES.r7.t0.t0.s4.clk )
    begin
        case ( \AES.r7.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t0.out  = { \AES.r7.t0.t0.k0 , \AES.r7.t0.t0.k0 , ( \AES.r7.t0.t0.k0  ^ \AES.r7.t0.t0.k1  ), \AES.r7.t0.t0.k1  };
    assign \AES.r7.t0.t1.clk  = \AES.r7.t0.clk ;
    assign \AES.r7.t0.t1.in  = \AES.r7.t0.b1 ;
    assign \AES.r7.t0.k1  = \AES.r7.t0.t1.out ;
    assign \AES.r7.t0.t1.s0.clk  = \AES.r7.t0.t1.clk ;
    assign \AES.r7.t0.t1.s0.in  = \AES.r7.t0.t1.in ;
    assign \AES.r7.t0.t1.k0  = \AES.r7.t0.t1.s0.out ;
    always @ (  posedge \AES.r7.t0.t1.s0.clk )
    begin
        case ( \AES.r7.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t1.s4.clk  = \AES.r7.t0.t1.clk ;
    assign \AES.r7.t0.t1.s4.in  = \AES.r7.t0.t1.in ;
    assign \AES.r7.t0.t1.k1  = \AES.r7.t0.t1.s4.out ;
    always @ (  posedge \AES.r7.t0.t1.s4.clk )
    begin
        case ( \AES.r7.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t1.out  = { \AES.r7.t0.t1.k0 , \AES.r7.t0.t1.k0 , ( \AES.r7.t0.t1.k0  ^ \AES.r7.t0.t1.k1  ), \AES.r7.t0.t1.k1  };
    assign \AES.r7.t0.t2.clk  = \AES.r7.t0.clk ;
    assign \AES.r7.t0.t2.in  = \AES.r7.t0.b2 ;
    assign \AES.r7.t0.k2  = \AES.r7.t0.t2.out ;
    assign \AES.r7.t0.t2.s0.clk  = \AES.r7.t0.t2.clk ;
    assign \AES.r7.t0.t2.s0.in  = \AES.r7.t0.t2.in ;
    assign \AES.r7.t0.t2.k0  = \AES.r7.t0.t2.s0.out ;
    always @ (  posedge \AES.r7.t0.t2.s0.clk )
    begin
        case ( \AES.r7.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t2.s4.clk  = \AES.r7.t0.t2.clk ;
    assign \AES.r7.t0.t2.s4.in  = \AES.r7.t0.t2.in ;
    assign \AES.r7.t0.t2.k1  = \AES.r7.t0.t2.s4.out ;
    always @ (  posedge \AES.r7.t0.t2.s4.clk )
    begin
        case ( \AES.r7.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t2.out  = { \AES.r7.t0.t2.k0 , \AES.r7.t0.t2.k0 , ( \AES.r7.t0.t2.k0  ^ \AES.r7.t0.t2.k1  ), \AES.r7.t0.t2.k1  };
    assign \AES.r7.t0.t3.clk  = \AES.r7.t0.clk ;
    assign \AES.r7.t0.t3.in  = \AES.r7.t0.b3 ;
    assign \AES.r7.t0.p3  = \AES.r7.t0.t3.out ;
    assign \AES.r7.t0.t3.s0.clk  = \AES.r7.t0.t3.clk ;
    assign \AES.r7.t0.t3.s0.in  = \AES.r7.t0.t3.in ;
    assign \AES.r7.t0.t3.k0  = \AES.r7.t0.t3.s0.out ;
    always @ (  posedge \AES.r7.t0.t3.s0.clk )
    begin
        case ( \AES.r7.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t3.s4.clk  = \AES.r7.t0.t3.clk ;
    assign \AES.r7.t0.t3.s4.in  = \AES.r7.t0.t3.in ;
    assign \AES.r7.t0.t3.k1  = \AES.r7.t0.t3.s4.out ;
    always @ (  posedge \AES.r7.t0.t3.s4.clk )
    begin
        case ( \AES.r7.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t0.t3.out  = { \AES.r7.t0.t3.k0 , \AES.r7.t0.t3.k0 , ( \AES.r7.t0.t3.k0  ^ \AES.r7.t0.t3.k1  ), \AES.r7.t0.t3.k1  };
    assign \AES.r7.t1.clk  = \AES.r7.clk ;
    assign \AES.r7.t1.state  = \AES.r7.s1 ;
    assign \AES.r7.p10  = \AES.r7.t1.p0 ;
    assign \AES.r7.p11  = \AES.r7.t1.p1 ;
    assign \AES.r7.p12  = \AES.r7.t1.p2 ;
    assign \AES.r7.p13  = \AES.r7.t1.p3 ;
    assign \AES.r7.t1.p0  = { \AES.r7.t1.k0 [7:0], \AES.r7.t1.k0 [31:8] };
    assign \AES.r7.t1.p1  = { \AES.r7.t1.k1 [15:0], \AES.r7.t1.k1 [31:16] };
    assign \AES.r7.t1.p2  = { \AES.r7.t1.k2 [23:0], \AES.r7.t1.k2 [31:24] };
    assign \AES.r7.t1.b0  = \AES.r7.t1.state [31:24];
    assign \AES.r7.t1.b1  = \AES.r7.t1.state [23:16];
    assign \AES.r7.t1.b2  = \AES.r7.t1.state [15:8];
    assign \AES.r7.t1.b3  = \AES.r7.t1.state [7:0];
    assign \AES.r7.t1.t0.clk  = \AES.r7.t1.clk ;
    assign \AES.r7.t1.t0.in  = \AES.r7.t1.b0 ;
    assign \AES.r7.t1.k0  = \AES.r7.t1.t0.out ;
    assign \AES.r7.t1.t0.s0.clk  = \AES.r7.t1.t0.clk ;
    assign \AES.r7.t1.t0.s0.in  = \AES.r7.t1.t0.in ;
    assign \AES.r7.t1.t0.k0  = \AES.r7.t1.t0.s0.out ;
    always @ (  posedge \AES.r7.t1.t0.s0.clk )
    begin
        case ( \AES.r7.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t0.s4.clk  = \AES.r7.t1.t0.clk ;
    assign \AES.r7.t1.t0.s4.in  = \AES.r7.t1.t0.in ;
    assign \AES.r7.t1.t0.k1  = \AES.r7.t1.t0.s4.out ;
    always @ (  posedge \AES.r7.t1.t0.s4.clk )
    begin
        case ( \AES.r7.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t0.out  = { \AES.r7.t1.t0.k0 , \AES.r7.t1.t0.k0 , ( \AES.r7.t1.t0.k0  ^ \AES.r7.t1.t0.k1  ), \AES.r7.t1.t0.k1  };
    assign \AES.r7.t1.t1.clk  = \AES.r7.t1.clk ;
    assign \AES.r7.t1.t1.in  = \AES.r7.t1.b1 ;
    assign \AES.r7.t1.k1  = \AES.r7.t1.t1.out ;
    assign \AES.r7.t1.t1.s0.clk  = \AES.r7.t1.t1.clk ;
    assign \AES.r7.t1.t1.s0.in  = \AES.r7.t1.t1.in ;
    assign \AES.r7.t1.t1.k0  = \AES.r7.t1.t1.s0.out ;
    always @ (  posedge \AES.r7.t1.t1.s0.clk )
    begin
        case ( \AES.r7.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t1.s4.clk  = \AES.r7.t1.t1.clk ;
    assign \AES.r7.t1.t1.s4.in  = \AES.r7.t1.t1.in ;
    assign \AES.r7.t1.t1.k1  = \AES.r7.t1.t1.s4.out ;
    always @ (  posedge \AES.r7.t1.t1.s4.clk )
    begin
        case ( \AES.r7.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t1.out  = { \AES.r7.t1.t1.k0 , \AES.r7.t1.t1.k0 , ( \AES.r7.t1.t1.k0  ^ \AES.r7.t1.t1.k1  ), \AES.r7.t1.t1.k1  };
    assign \AES.r7.t1.t2.clk  = \AES.r7.t1.clk ;
    assign \AES.r7.t1.t2.in  = \AES.r7.t1.b2 ;
    assign \AES.r7.t1.k2  = \AES.r7.t1.t2.out ;
    assign \AES.r7.t1.t2.s0.clk  = \AES.r7.t1.t2.clk ;
    assign \AES.r7.t1.t2.s0.in  = \AES.r7.t1.t2.in ;
    assign \AES.r7.t1.t2.k0  = \AES.r7.t1.t2.s0.out ;
    always @ (  posedge \AES.r7.t1.t2.s0.clk )
    begin
        case ( \AES.r7.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t2.s4.clk  = \AES.r7.t1.t2.clk ;
    assign \AES.r7.t1.t2.s4.in  = \AES.r7.t1.t2.in ;
    assign \AES.r7.t1.t2.k1  = \AES.r7.t1.t2.s4.out ;
    always @ (  posedge \AES.r7.t1.t2.s4.clk )
    begin
        case ( \AES.r7.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t2.out  = { \AES.r7.t1.t2.k0 , \AES.r7.t1.t2.k0 , ( \AES.r7.t1.t2.k0  ^ \AES.r7.t1.t2.k1  ), \AES.r7.t1.t2.k1  };
    assign \AES.r7.t1.t3.clk  = \AES.r7.t1.clk ;
    assign \AES.r7.t1.t3.in  = \AES.r7.t1.b3 ;
    assign \AES.r7.t1.p3  = \AES.r7.t1.t3.out ;
    assign \AES.r7.t1.t3.s0.clk  = \AES.r7.t1.t3.clk ;
    assign \AES.r7.t1.t3.s0.in  = \AES.r7.t1.t3.in ;
    assign \AES.r7.t1.t3.k0  = \AES.r7.t1.t3.s0.out ;
    always @ (  posedge \AES.r7.t1.t3.s0.clk )
    begin
        case ( \AES.r7.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t3.s4.clk  = \AES.r7.t1.t3.clk ;
    assign \AES.r7.t1.t3.s4.in  = \AES.r7.t1.t3.in ;
    assign \AES.r7.t1.t3.k1  = \AES.r7.t1.t3.s4.out ;
    always @ (  posedge \AES.r7.t1.t3.s4.clk )
    begin
        case ( \AES.r7.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t1.t3.out  = { \AES.r7.t1.t3.k0 , \AES.r7.t1.t3.k0 , ( \AES.r7.t1.t3.k0  ^ \AES.r7.t1.t3.k1  ), \AES.r7.t1.t3.k1  };
    assign \AES.r7.t2.clk  = \AES.r7.clk ;
    assign \AES.r7.t2.state  = \AES.r7.s2 ;
    assign \AES.r7.p20  = \AES.r7.t2.p0 ;
    assign \AES.r7.p21  = \AES.r7.t2.p1 ;
    assign \AES.r7.p22  = \AES.r7.t2.p2 ;
    assign \AES.r7.p23  = \AES.r7.t2.p3 ;
    assign \AES.r7.t2.p0  = { \AES.r7.t2.k0 [7:0], \AES.r7.t2.k0 [31:8] };
    assign \AES.r7.t2.p1  = { \AES.r7.t2.k1 [15:0], \AES.r7.t2.k1 [31:16] };
    assign \AES.r7.t2.p2  = { \AES.r7.t2.k2 [23:0], \AES.r7.t2.k2 [31:24] };
    assign \AES.r7.t2.b0  = \AES.r7.t2.state [31:24];
    assign \AES.r7.t2.b1  = \AES.r7.t2.state [23:16];
    assign \AES.r7.t2.b2  = \AES.r7.t2.state [15:8];
    assign \AES.r7.t2.b3  = \AES.r7.t2.state [7:0];
    assign \AES.r7.t2.t0.clk  = \AES.r7.t2.clk ;
    assign \AES.r7.t2.t0.in  = \AES.r7.t2.b0 ;
    assign \AES.r7.t2.k0  = \AES.r7.t2.t0.out ;
    assign \AES.r7.t2.t0.s0.clk  = \AES.r7.t2.t0.clk ;
    assign \AES.r7.t2.t0.s0.in  = \AES.r7.t2.t0.in ;
    assign \AES.r7.t2.t0.k0  = \AES.r7.t2.t0.s0.out ;
    always @ (  posedge \AES.r7.t2.t0.s0.clk )
    begin
        case ( \AES.r7.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t0.s4.clk  = \AES.r7.t2.t0.clk ;
    assign \AES.r7.t2.t0.s4.in  = \AES.r7.t2.t0.in ;
    assign \AES.r7.t2.t0.k1  = \AES.r7.t2.t0.s4.out ;
    always @ (  posedge \AES.r7.t2.t0.s4.clk )
    begin
        case ( \AES.r7.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t0.out  = { \AES.r7.t2.t0.k0 , \AES.r7.t2.t0.k0 , ( \AES.r7.t2.t0.k0  ^ \AES.r7.t2.t0.k1  ), \AES.r7.t2.t0.k1  };
    assign \AES.r7.t2.t1.clk  = \AES.r7.t2.clk ;
    assign \AES.r7.t2.t1.in  = \AES.r7.t2.b1 ;
    assign \AES.r7.t2.k1  = \AES.r7.t2.t1.out ;
    assign \AES.r7.t2.t1.s0.clk  = \AES.r7.t2.t1.clk ;
    assign \AES.r7.t2.t1.s0.in  = \AES.r7.t2.t1.in ;
    assign \AES.r7.t2.t1.k0  = \AES.r7.t2.t1.s0.out ;
    always @ (  posedge \AES.r7.t2.t1.s0.clk )
    begin
        case ( \AES.r7.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t1.s4.clk  = \AES.r7.t2.t1.clk ;
    assign \AES.r7.t2.t1.s4.in  = \AES.r7.t2.t1.in ;
    assign \AES.r7.t2.t1.k1  = \AES.r7.t2.t1.s4.out ;
    always @ (  posedge \AES.r7.t2.t1.s4.clk )
    begin
        case ( \AES.r7.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t1.out  = { \AES.r7.t2.t1.k0 , \AES.r7.t2.t1.k0 , ( \AES.r7.t2.t1.k0  ^ \AES.r7.t2.t1.k1  ), \AES.r7.t2.t1.k1  };
    assign \AES.r7.t2.t2.clk  = \AES.r7.t2.clk ;
    assign \AES.r7.t2.t2.in  = \AES.r7.t2.b2 ;
    assign \AES.r7.t2.k2  = \AES.r7.t2.t2.out ;
    assign \AES.r7.t2.t2.s0.clk  = \AES.r7.t2.t2.clk ;
    assign \AES.r7.t2.t2.s0.in  = \AES.r7.t2.t2.in ;
    assign \AES.r7.t2.t2.k0  = \AES.r7.t2.t2.s0.out ;
    always @ (  posedge \AES.r7.t2.t2.s0.clk )
    begin
        case ( \AES.r7.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t2.s4.clk  = \AES.r7.t2.t2.clk ;
    assign \AES.r7.t2.t2.s4.in  = \AES.r7.t2.t2.in ;
    assign \AES.r7.t2.t2.k1  = \AES.r7.t2.t2.s4.out ;
    always @ (  posedge \AES.r7.t2.t2.s4.clk )
    begin
        case ( \AES.r7.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t2.out  = { \AES.r7.t2.t2.k0 , \AES.r7.t2.t2.k0 , ( \AES.r7.t2.t2.k0  ^ \AES.r7.t2.t2.k1  ), \AES.r7.t2.t2.k1  };
    assign \AES.r7.t2.t3.clk  = \AES.r7.t2.clk ;
    assign \AES.r7.t2.t3.in  = \AES.r7.t2.b3 ;
    assign \AES.r7.t2.p3  = \AES.r7.t2.t3.out ;
    assign \AES.r7.t2.t3.s0.clk  = \AES.r7.t2.t3.clk ;
    assign \AES.r7.t2.t3.s0.in  = \AES.r7.t2.t3.in ;
    assign \AES.r7.t2.t3.k0  = \AES.r7.t2.t3.s0.out ;
    always @ (  posedge \AES.r7.t2.t3.s0.clk )
    begin
        case ( \AES.r7.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t3.s4.clk  = \AES.r7.t2.t3.clk ;
    assign \AES.r7.t2.t3.s4.in  = \AES.r7.t2.t3.in ;
    assign \AES.r7.t2.t3.k1  = \AES.r7.t2.t3.s4.out ;
    always @ (  posedge \AES.r7.t2.t3.s4.clk )
    begin
        case ( \AES.r7.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t2.t3.out  = { \AES.r7.t2.t3.k0 , \AES.r7.t2.t3.k0 , ( \AES.r7.t2.t3.k0  ^ \AES.r7.t2.t3.k1  ), \AES.r7.t2.t3.k1  };
    assign \AES.r7.t3.clk  = \AES.r7.clk ;
    assign \AES.r7.t3.state  = \AES.r7.s3 ;
    assign \AES.r7.p30  = \AES.r7.t3.p0 ;
    assign \AES.r7.p31  = \AES.r7.t3.p1 ;
    assign \AES.r7.p32  = \AES.r7.t3.p2 ;
    assign \AES.r7.p33  = \AES.r7.t3.p3 ;
    assign \AES.r7.t3.p0  = { \AES.r7.t3.k0 [7:0], \AES.r7.t3.k0 [31:8] };
    assign \AES.r7.t3.p1  = { \AES.r7.t3.k1 [15:0], \AES.r7.t3.k1 [31:16] };
    assign \AES.r7.t3.p2  = { \AES.r7.t3.k2 [23:0], \AES.r7.t3.k2 [31:24] };
    assign \AES.r7.t3.b0  = \AES.r7.t3.state [31:24];
    assign \AES.r7.t3.b1  = \AES.r7.t3.state [23:16];
    assign \AES.r7.t3.b2  = \AES.r7.t3.state [15:8];
    assign \AES.r7.t3.b3  = \AES.r7.t3.state [7:0];
    assign \AES.r7.t3.t0.clk  = \AES.r7.t3.clk ;
    assign \AES.r7.t3.t0.in  = \AES.r7.t3.b0 ;
    assign \AES.r7.t3.k0  = \AES.r7.t3.t0.out ;
    assign \AES.r7.t3.t0.s0.clk  = \AES.r7.t3.t0.clk ;
    assign \AES.r7.t3.t0.s0.in  = \AES.r7.t3.t0.in ;
    assign \AES.r7.t3.t0.k0  = \AES.r7.t3.t0.s0.out ;
    always @ (  posedge \AES.r7.t3.t0.s0.clk )
    begin
        case ( \AES.r7.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t0.s4.clk  = \AES.r7.t3.t0.clk ;
    assign \AES.r7.t3.t0.s4.in  = \AES.r7.t3.t0.in ;
    assign \AES.r7.t3.t0.k1  = \AES.r7.t3.t0.s4.out ;
    always @ (  posedge \AES.r7.t3.t0.s4.clk )
    begin
        case ( \AES.r7.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t0.out  = { \AES.r7.t3.t0.k0 , \AES.r7.t3.t0.k0 , ( \AES.r7.t3.t0.k0  ^ \AES.r7.t3.t0.k1  ), \AES.r7.t3.t0.k1  };
    assign \AES.r7.t3.t1.clk  = \AES.r7.t3.clk ;
    assign \AES.r7.t3.t1.in  = \AES.r7.t3.b1 ;
    assign \AES.r7.t3.k1  = \AES.r7.t3.t1.out ;
    assign \AES.r7.t3.t1.s0.clk  = \AES.r7.t3.t1.clk ;
    assign \AES.r7.t3.t1.s0.in  = \AES.r7.t3.t1.in ;
    assign \AES.r7.t3.t1.k0  = \AES.r7.t3.t1.s0.out ;
    always @ (  posedge \AES.r7.t3.t1.s0.clk )
    begin
        case ( \AES.r7.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t1.s4.clk  = \AES.r7.t3.t1.clk ;
    assign \AES.r7.t3.t1.s4.in  = \AES.r7.t3.t1.in ;
    assign \AES.r7.t3.t1.k1  = \AES.r7.t3.t1.s4.out ;
    always @ (  posedge \AES.r7.t3.t1.s4.clk )
    begin
        case ( \AES.r7.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t1.out  = { \AES.r7.t3.t1.k0 , \AES.r7.t3.t1.k0 , ( \AES.r7.t3.t1.k0  ^ \AES.r7.t3.t1.k1  ), \AES.r7.t3.t1.k1  };
    assign \AES.r7.t3.t2.clk  = \AES.r7.t3.clk ;
    assign \AES.r7.t3.t2.in  = \AES.r7.t3.b2 ;
    assign \AES.r7.t3.k2  = \AES.r7.t3.t2.out ;
    assign \AES.r7.t3.t2.s0.clk  = \AES.r7.t3.t2.clk ;
    assign \AES.r7.t3.t2.s0.in  = \AES.r7.t3.t2.in ;
    assign \AES.r7.t3.t2.k0  = \AES.r7.t3.t2.s0.out ;
    always @ (  posedge \AES.r7.t3.t2.s0.clk )
    begin
        case ( \AES.r7.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t2.s4.clk  = \AES.r7.t3.t2.clk ;
    assign \AES.r7.t3.t2.s4.in  = \AES.r7.t3.t2.in ;
    assign \AES.r7.t3.t2.k1  = \AES.r7.t3.t2.s4.out ;
    always @ (  posedge \AES.r7.t3.t2.s4.clk )
    begin
        case ( \AES.r7.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t2.out  = { \AES.r7.t3.t2.k0 , \AES.r7.t3.t2.k0 , ( \AES.r7.t3.t2.k0  ^ \AES.r7.t3.t2.k1  ), \AES.r7.t3.t2.k1  };
    assign \AES.r7.t3.t3.clk  = \AES.r7.t3.clk ;
    assign \AES.r7.t3.t3.in  = \AES.r7.t3.b3 ;
    assign \AES.r7.t3.p3  = \AES.r7.t3.t3.out ;
    assign \AES.r7.t3.t3.s0.clk  = \AES.r7.t3.t3.clk ;
    assign \AES.r7.t3.t3.s0.in  = \AES.r7.t3.t3.in ;
    assign \AES.r7.t3.t3.k0  = \AES.r7.t3.t3.s0.out ;
    always @ (  posedge \AES.r7.t3.t3.s0.clk )
    begin
        case ( \AES.r7.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t3.s4.clk  = \AES.r7.t3.t3.clk ;
    assign \AES.r7.t3.t3.s4.in  = \AES.r7.t3.t3.in ;
    assign \AES.r7.t3.t3.k1  = \AES.r7.t3.t3.s4.out ;
    always @ (  posedge \AES.r7.t3.t3.s4.clk )
    begin
        case ( \AES.r7.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r7.t3.t3.out  = { \AES.r7.t3.t3.k0 , \AES.r7.t3.t3.k0 , ( \AES.r7.t3.t3.k0  ^ \AES.r7.t3.t3.k1  ), \AES.r7.t3.t3.k1  };
    assign \AES.r7.z0  = ( ( ( ( \AES.r7.p00  ^ \AES.r7.p11  ) ^ \AES.r7.p22  ) ^ \AES.r7.p33  ) ^ \AES.r7.k0  );
    assign \AES.r7.z1  = ( ( ( ( \AES.r7.p03  ^ \AES.r7.p10  ) ^ \AES.r7.p21  ) ^ \AES.r7.p32  ) ^ \AES.r7.k1  );
    assign \AES.r7.z2  = ( ( ( ( \AES.r7.p02  ^ \AES.r7.p13  ) ^ \AES.r7.p20  ) ^ \AES.r7.p31  ) ^ \AES.r7.k2  );
    assign \AES.r7.z3  = ( ( ( ( \AES.r7.p01  ^ \AES.r7.p12  ) ^ \AES.r7.p23  ) ^ \AES.r7.p30  ) ^ \AES.r7.k3  );
    always @ (  posedge \AES.r7.clk )
    begin
    end
    assign \AES.r8.clk  = \AES.clk ;
    assign \AES.r8.state_in  = \AES.s7 ;
    assign \AES.r8.key  = \AES.k7b ;
    assign \AES.s8  = \AES.r8.state_out ;
    assign \AES.r8.k0  = \AES.r8.key [127:96];
    assign \AES.r8.k1  = \AES.r8.key [95:64];
    assign \AES.r8.k2  = \AES.r8.key [63:32];
    assign \AES.r8.k3  = \AES.r8.key [31:0];
    assign \AES.r8.s0  = \AES.r8.state_in [127:96];
    assign \AES.r8.s1  = \AES.r8.state_in [95:64];
    assign \AES.r8.s2  = \AES.r8.state_in [63:32];
    assign \AES.r8.s3  = \AES.r8.state_in [31:0];
    assign \AES.r8.t0.clk  = \AES.r8.clk ;
    assign \AES.r8.t0.state  = \AES.r8.s0 ;
    assign \AES.r8.p00  = \AES.r8.t0.p0 ;
    assign \AES.r8.p01  = \AES.r8.t0.p1 ;
    assign \AES.r8.p02  = \AES.r8.t0.p2 ;
    assign \AES.r8.p03  = \AES.r8.t0.p3 ;
    assign \AES.r8.t0.p0  = { \AES.r8.t0.k0 [7:0], \AES.r8.t0.k0 [31:8] };
    assign \AES.r8.t0.p1  = { \AES.r8.t0.k1 [15:0], \AES.r8.t0.k1 [31:16] };
    assign \AES.r8.t0.p2  = { \AES.r8.t0.k2 [23:0], \AES.r8.t0.k2 [31:24] };
    assign \AES.r8.t0.b0  = \AES.r8.t0.state [31:24];
    assign \AES.r8.t0.b1  = \AES.r8.t0.state [23:16];
    assign \AES.r8.t0.b2  = \AES.r8.t0.state [15:8];
    assign \AES.r8.t0.b3  = \AES.r8.t0.state [7:0];
    assign \AES.r8.t0.t0.clk  = \AES.r8.t0.clk ;
    assign \AES.r8.t0.t0.in  = \AES.r8.t0.b0 ;
    assign \AES.r8.t0.k0  = \AES.r8.t0.t0.out ;
    assign \AES.r8.t0.t0.s0.clk  = \AES.r8.t0.t0.clk ;
    assign \AES.r8.t0.t0.s0.in  = \AES.r8.t0.t0.in ;
    assign \AES.r8.t0.t0.k0  = \AES.r8.t0.t0.s0.out ;
    always @ (  posedge \AES.r8.t0.t0.s0.clk )
    begin
        case ( \AES.r8.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t0.s4.clk  = \AES.r8.t0.t0.clk ;
    assign \AES.r8.t0.t0.s4.in  = \AES.r8.t0.t0.in ;
    assign \AES.r8.t0.t0.k1  = \AES.r8.t0.t0.s4.out ;
    always @ (  posedge \AES.r8.t0.t0.s4.clk )
    begin
        case ( \AES.r8.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t0.out  = { \AES.r8.t0.t0.k0 , \AES.r8.t0.t0.k0 , ( \AES.r8.t0.t0.k0  ^ \AES.r8.t0.t0.k1  ), \AES.r8.t0.t0.k1  };
    assign \AES.r8.t0.t1.clk  = \AES.r8.t0.clk ;
    assign \AES.r8.t0.t1.in  = \AES.r8.t0.b1 ;
    assign \AES.r8.t0.k1  = \AES.r8.t0.t1.out ;
    assign \AES.r8.t0.t1.s0.clk  = \AES.r8.t0.t1.clk ;
    assign \AES.r8.t0.t1.s0.in  = \AES.r8.t0.t1.in ;
    assign \AES.r8.t0.t1.k0  = \AES.r8.t0.t1.s0.out ;
    always @ (  posedge \AES.r8.t0.t1.s0.clk )
    begin
        case ( \AES.r8.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t1.s4.clk  = \AES.r8.t0.t1.clk ;
    assign \AES.r8.t0.t1.s4.in  = \AES.r8.t0.t1.in ;
    assign \AES.r8.t0.t1.k1  = \AES.r8.t0.t1.s4.out ;
    always @ (  posedge \AES.r8.t0.t1.s4.clk )
    begin
        case ( \AES.r8.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t1.out  = { \AES.r8.t0.t1.k0 , \AES.r8.t0.t1.k0 , ( \AES.r8.t0.t1.k0  ^ \AES.r8.t0.t1.k1  ), \AES.r8.t0.t1.k1  };
    assign \AES.r8.t0.t2.clk  = \AES.r8.t0.clk ;
    assign \AES.r8.t0.t2.in  = \AES.r8.t0.b2 ;
    assign \AES.r8.t0.k2  = \AES.r8.t0.t2.out ;
    assign \AES.r8.t0.t2.s0.clk  = \AES.r8.t0.t2.clk ;
    assign \AES.r8.t0.t2.s0.in  = \AES.r8.t0.t2.in ;
    assign \AES.r8.t0.t2.k0  = \AES.r8.t0.t2.s0.out ;
    always @ (  posedge \AES.r8.t0.t2.s0.clk )
    begin
        case ( \AES.r8.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t2.s4.clk  = \AES.r8.t0.t2.clk ;
    assign \AES.r8.t0.t2.s4.in  = \AES.r8.t0.t2.in ;
    assign \AES.r8.t0.t2.k1  = \AES.r8.t0.t2.s4.out ;
    always @ (  posedge \AES.r8.t0.t2.s4.clk )
    begin
        case ( \AES.r8.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t2.out  = { \AES.r8.t0.t2.k0 , \AES.r8.t0.t2.k0 , ( \AES.r8.t0.t2.k0  ^ \AES.r8.t0.t2.k1  ), \AES.r8.t0.t2.k1  };
    assign \AES.r8.t0.t3.clk  = \AES.r8.t0.clk ;
    assign \AES.r8.t0.t3.in  = \AES.r8.t0.b3 ;
    assign \AES.r8.t0.p3  = \AES.r8.t0.t3.out ;
    assign \AES.r8.t0.t3.s0.clk  = \AES.r8.t0.t3.clk ;
    assign \AES.r8.t0.t3.s0.in  = \AES.r8.t0.t3.in ;
    assign \AES.r8.t0.t3.k0  = \AES.r8.t0.t3.s0.out ;
    always @ (  posedge \AES.r8.t0.t3.s0.clk )
    begin
        case ( \AES.r8.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t3.s4.clk  = \AES.r8.t0.t3.clk ;
    assign \AES.r8.t0.t3.s4.in  = \AES.r8.t0.t3.in ;
    assign \AES.r8.t0.t3.k1  = \AES.r8.t0.t3.s4.out ;
    always @ (  posedge \AES.r8.t0.t3.s4.clk )
    begin
        case ( \AES.r8.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t0.t3.out  = { \AES.r8.t0.t3.k0 , \AES.r8.t0.t3.k0 , ( \AES.r8.t0.t3.k0  ^ \AES.r8.t0.t3.k1  ), \AES.r8.t0.t3.k1  };
    assign \AES.r8.t1.clk  = \AES.r8.clk ;
    assign \AES.r8.t1.state  = \AES.r8.s1 ;
    assign \AES.r8.p10  = \AES.r8.t1.p0 ;
    assign \AES.r8.p11  = \AES.r8.t1.p1 ;
    assign \AES.r8.p12  = \AES.r8.t1.p2 ;
    assign \AES.r8.p13  = \AES.r8.t1.p3 ;
    assign \AES.r8.t1.p0  = { \AES.r8.t1.k0 [7:0], \AES.r8.t1.k0 [31:8] };
    assign \AES.r8.t1.p1  = { \AES.r8.t1.k1 [15:0], \AES.r8.t1.k1 [31:16] };
    assign \AES.r8.t1.p2  = { \AES.r8.t1.k2 [23:0], \AES.r8.t1.k2 [31:24] };
    assign \AES.r8.t1.b0  = \AES.r8.t1.state [31:24];
    assign \AES.r8.t1.b1  = \AES.r8.t1.state [23:16];
    assign \AES.r8.t1.b2  = \AES.r8.t1.state [15:8];
    assign \AES.r8.t1.b3  = \AES.r8.t1.state [7:0];
    assign \AES.r8.t1.t0.clk  = \AES.r8.t1.clk ;
    assign \AES.r8.t1.t0.in  = \AES.r8.t1.b0 ;
    assign \AES.r8.t1.k0  = \AES.r8.t1.t0.out ;
    assign \AES.r8.t1.t0.s0.clk  = \AES.r8.t1.t0.clk ;
    assign \AES.r8.t1.t0.s0.in  = \AES.r8.t1.t0.in ;
    assign \AES.r8.t1.t0.k0  = \AES.r8.t1.t0.s0.out ;
    always @ (  posedge \AES.r8.t1.t0.s0.clk )
    begin
        case ( \AES.r8.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t0.s4.clk  = \AES.r8.t1.t0.clk ;
    assign \AES.r8.t1.t0.s4.in  = \AES.r8.t1.t0.in ;
    assign \AES.r8.t1.t0.k1  = \AES.r8.t1.t0.s4.out ;
    always @ (  posedge \AES.r8.t1.t0.s4.clk )
    begin
        case ( \AES.r8.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t0.out  = { \AES.r8.t1.t0.k0 , \AES.r8.t1.t0.k0 , ( \AES.r8.t1.t0.k0  ^ \AES.r8.t1.t0.k1  ), \AES.r8.t1.t0.k1  };
    assign \AES.r8.t1.t1.clk  = \AES.r8.t1.clk ;
    assign \AES.r8.t1.t1.in  = \AES.r8.t1.b1 ;
    assign \AES.r8.t1.k1  = \AES.r8.t1.t1.out ;
    assign \AES.r8.t1.t1.s0.clk  = \AES.r8.t1.t1.clk ;
    assign \AES.r8.t1.t1.s0.in  = \AES.r8.t1.t1.in ;
    assign \AES.r8.t1.t1.k0  = \AES.r8.t1.t1.s0.out ;
    always @ (  posedge \AES.r8.t1.t1.s0.clk )
    begin
        case ( \AES.r8.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t1.s4.clk  = \AES.r8.t1.t1.clk ;
    assign \AES.r8.t1.t1.s4.in  = \AES.r8.t1.t1.in ;
    assign \AES.r8.t1.t1.k1  = \AES.r8.t1.t1.s4.out ;
    always @ (  posedge \AES.r8.t1.t1.s4.clk )
    begin
        case ( \AES.r8.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t1.out  = { \AES.r8.t1.t1.k0 , \AES.r8.t1.t1.k0 , ( \AES.r8.t1.t1.k0  ^ \AES.r8.t1.t1.k1  ), \AES.r8.t1.t1.k1  };
    assign \AES.r8.t1.t2.clk  = \AES.r8.t1.clk ;
    assign \AES.r8.t1.t2.in  = \AES.r8.t1.b2 ;
    assign \AES.r8.t1.k2  = \AES.r8.t1.t2.out ;
    assign \AES.r8.t1.t2.s0.clk  = \AES.r8.t1.t2.clk ;
    assign \AES.r8.t1.t2.s0.in  = \AES.r8.t1.t2.in ;
    assign \AES.r8.t1.t2.k0  = \AES.r8.t1.t2.s0.out ;
    always @ (  posedge \AES.r8.t1.t2.s0.clk )
    begin
        case ( \AES.r8.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t2.s4.clk  = \AES.r8.t1.t2.clk ;
    assign \AES.r8.t1.t2.s4.in  = \AES.r8.t1.t2.in ;
    assign \AES.r8.t1.t2.k1  = \AES.r8.t1.t2.s4.out ;
    always @ (  posedge \AES.r8.t1.t2.s4.clk )
    begin
        case ( \AES.r8.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t2.out  = { \AES.r8.t1.t2.k0 , \AES.r8.t1.t2.k0 , ( \AES.r8.t1.t2.k0  ^ \AES.r8.t1.t2.k1  ), \AES.r8.t1.t2.k1  };
    assign \AES.r8.t1.t3.clk  = \AES.r8.t1.clk ;
    assign \AES.r8.t1.t3.in  = \AES.r8.t1.b3 ;
    assign \AES.r8.t1.p3  = \AES.r8.t1.t3.out ;
    assign \AES.r8.t1.t3.s0.clk  = \AES.r8.t1.t3.clk ;
    assign \AES.r8.t1.t3.s0.in  = \AES.r8.t1.t3.in ;
    assign \AES.r8.t1.t3.k0  = \AES.r8.t1.t3.s0.out ;
    always @ (  posedge \AES.r8.t1.t3.s0.clk )
    begin
        case ( \AES.r8.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t3.s4.clk  = \AES.r8.t1.t3.clk ;
    assign \AES.r8.t1.t3.s4.in  = \AES.r8.t1.t3.in ;
    assign \AES.r8.t1.t3.k1  = \AES.r8.t1.t3.s4.out ;
    always @ (  posedge \AES.r8.t1.t3.s4.clk )
    begin
        case ( \AES.r8.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t1.t3.out  = { \AES.r8.t1.t3.k0 , \AES.r8.t1.t3.k0 , ( \AES.r8.t1.t3.k0  ^ \AES.r8.t1.t3.k1  ), \AES.r8.t1.t3.k1  };
    assign \AES.r8.t2.clk  = \AES.r8.clk ;
    assign \AES.r8.t2.state  = \AES.r8.s2 ;
    assign \AES.r8.p20  = \AES.r8.t2.p0 ;
    assign \AES.r8.p21  = \AES.r8.t2.p1 ;
    assign \AES.r8.p22  = \AES.r8.t2.p2 ;
    assign \AES.r8.p23  = \AES.r8.t2.p3 ;
    assign \AES.r8.t2.p0  = { \AES.r8.t2.k0 [7:0], \AES.r8.t2.k0 [31:8] };
    assign \AES.r8.t2.p1  = { \AES.r8.t2.k1 [15:0], \AES.r8.t2.k1 [31:16] };
    assign \AES.r8.t2.p2  = { \AES.r8.t2.k2 [23:0], \AES.r8.t2.k2 [31:24] };
    assign \AES.r8.t2.b0  = \AES.r8.t2.state [31:24];
    assign \AES.r8.t2.b1  = \AES.r8.t2.state [23:16];
    assign \AES.r8.t2.b2  = \AES.r8.t2.state [15:8];
    assign \AES.r8.t2.b3  = \AES.r8.t2.state [7:0];
    assign \AES.r8.t2.t0.clk  = \AES.r8.t2.clk ;
    assign \AES.r8.t2.t0.in  = \AES.r8.t2.b0 ;
    assign \AES.r8.t2.k0  = \AES.r8.t2.t0.out ;
    assign \AES.r8.t2.t0.s0.clk  = \AES.r8.t2.t0.clk ;
    assign \AES.r8.t2.t0.s0.in  = \AES.r8.t2.t0.in ;
    assign \AES.r8.t2.t0.k0  = \AES.r8.t2.t0.s0.out ;
    always @ (  posedge \AES.r8.t2.t0.s0.clk )
    begin
        case ( \AES.r8.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t0.s4.clk  = \AES.r8.t2.t0.clk ;
    assign \AES.r8.t2.t0.s4.in  = \AES.r8.t2.t0.in ;
    assign \AES.r8.t2.t0.k1  = \AES.r8.t2.t0.s4.out ;
    always @ (  posedge \AES.r8.t2.t0.s4.clk )
    begin
        case ( \AES.r8.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t0.out  = { \AES.r8.t2.t0.k0 , \AES.r8.t2.t0.k0 , ( \AES.r8.t2.t0.k0  ^ \AES.r8.t2.t0.k1  ), \AES.r8.t2.t0.k1  };
    assign \AES.r8.t2.t1.clk  = \AES.r8.t2.clk ;
    assign \AES.r8.t2.t1.in  = \AES.r8.t2.b1 ;
    assign \AES.r8.t2.k1  = \AES.r8.t2.t1.out ;
    assign \AES.r8.t2.t1.s0.clk  = \AES.r8.t2.t1.clk ;
    assign \AES.r8.t2.t1.s0.in  = \AES.r8.t2.t1.in ;
    assign \AES.r8.t2.t1.k0  = \AES.r8.t2.t1.s0.out ;
    always @ (  posedge \AES.r8.t2.t1.s0.clk )
    begin
        case ( \AES.r8.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t1.s4.clk  = \AES.r8.t2.t1.clk ;
    assign \AES.r8.t2.t1.s4.in  = \AES.r8.t2.t1.in ;
    assign \AES.r8.t2.t1.k1  = \AES.r8.t2.t1.s4.out ;
    always @ (  posedge \AES.r8.t2.t1.s4.clk )
    begin
        case ( \AES.r8.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t1.out  = { \AES.r8.t2.t1.k0 , \AES.r8.t2.t1.k0 , ( \AES.r8.t2.t1.k0  ^ \AES.r8.t2.t1.k1  ), \AES.r8.t2.t1.k1  };
    assign \AES.r8.t2.t2.clk  = \AES.r8.t2.clk ;
    assign \AES.r8.t2.t2.in  = \AES.r8.t2.b2 ;
    assign \AES.r8.t2.k2  = \AES.r8.t2.t2.out ;
    assign \AES.r8.t2.t2.s0.clk  = \AES.r8.t2.t2.clk ;
    assign \AES.r8.t2.t2.s0.in  = \AES.r8.t2.t2.in ;
    assign \AES.r8.t2.t2.k0  = \AES.r8.t2.t2.s0.out ;
    always @ (  posedge \AES.r8.t2.t2.s0.clk )
    begin
        case ( \AES.r8.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t2.s4.clk  = \AES.r8.t2.t2.clk ;
    assign \AES.r8.t2.t2.s4.in  = \AES.r8.t2.t2.in ;
    assign \AES.r8.t2.t2.k1  = \AES.r8.t2.t2.s4.out ;
    always @ (  posedge \AES.r8.t2.t2.s4.clk )
    begin
        case ( \AES.r8.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t2.out  = { \AES.r8.t2.t2.k0 , \AES.r8.t2.t2.k0 , ( \AES.r8.t2.t2.k0  ^ \AES.r8.t2.t2.k1  ), \AES.r8.t2.t2.k1  };
    assign \AES.r8.t2.t3.clk  = \AES.r8.t2.clk ;
    assign \AES.r8.t2.t3.in  = \AES.r8.t2.b3 ;
    assign \AES.r8.t2.p3  = \AES.r8.t2.t3.out ;
    assign \AES.r8.t2.t3.s0.clk  = \AES.r8.t2.t3.clk ;
    assign \AES.r8.t2.t3.s0.in  = \AES.r8.t2.t3.in ;
    assign \AES.r8.t2.t3.k0  = \AES.r8.t2.t3.s0.out ;
    always @ (  posedge \AES.r8.t2.t3.s0.clk )
    begin
        case ( \AES.r8.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t3.s4.clk  = \AES.r8.t2.t3.clk ;
    assign \AES.r8.t2.t3.s4.in  = \AES.r8.t2.t3.in ;
    assign \AES.r8.t2.t3.k1  = \AES.r8.t2.t3.s4.out ;
    always @ (  posedge \AES.r8.t2.t3.s4.clk )
    begin
        case ( \AES.r8.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t2.t3.out  = { \AES.r8.t2.t3.k0 , \AES.r8.t2.t3.k0 , ( \AES.r8.t2.t3.k0  ^ \AES.r8.t2.t3.k1  ), \AES.r8.t2.t3.k1  };
    assign \AES.r8.t3.clk  = \AES.r8.clk ;
    assign \AES.r8.t3.state  = \AES.r8.s3 ;
    assign \AES.r8.p30  = \AES.r8.t3.p0 ;
    assign \AES.r8.p31  = \AES.r8.t3.p1 ;
    assign \AES.r8.p32  = \AES.r8.t3.p2 ;
    assign \AES.r8.p33  = \AES.r8.t3.p3 ;
    assign \AES.r8.t3.p0  = { \AES.r8.t3.k0 [7:0], \AES.r8.t3.k0 [31:8] };
    assign \AES.r8.t3.p1  = { \AES.r8.t3.k1 [15:0], \AES.r8.t3.k1 [31:16] };
    assign \AES.r8.t3.p2  = { \AES.r8.t3.k2 [23:0], \AES.r8.t3.k2 [31:24] };
    assign \AES.r8.t3.b0  = \AES.r8.t3.state [31:24];
    assign \AES.r8.t3.b1  = \AES.r8.t3.state [23:16];
    assign \AES.r8.t3.b2  = \AES.r8.t3.state [15:8];
    assign \AES.r8.t3.b3  = \AES.r8.t3.state [7:0];
    assign \AES.r8.t3.t0.clk  = \AES.r8.t3.clk ;
    assign \AES.r8.t3.t0.in  = \AES.r8.t3.b0 ;
    assign \AES.r8.t3.k0  = \AES.r8.t3.t0.out ;
    assign \AES.r8.t3.t0.s0.clk  = \AES.r8.t3.t0.clk ;
    assign \AES.r8.t3.t0.s0.in  = \AES.r8.t3.t0.in ;
    assign \AES.r8.t3.t0.k0  = \AES.r8.t3.t0.s0.out ;
    always @ (  posedge \AES.r8.t3.t0.s0.clk )
    begin
        case ( \AES.r8.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t0.s4.clk  = \AES.r8.t3.t0.clk ;
    assign \AES.r8.t3.t0.s4.in  = \AES.r8.t3.t0.in ;
    assign \AES.r8.t3.t0.k1  = \AES.r8.t3.t0.s4.out ;
    always @ (  posedge \AES.r8.t3.t0.s4.clk )
    begin
        case ( \AES.r8.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t0.out  = { \AES.r8.t3.t0.k0 , \AES.r8.t3.t0.k0 , ( \AES.r8.t3.t0.k0  ^ \AES.r8.t3.t0.k1  ), \AES.r8.t3.t0.k1  };
    assign \AES.r8.t3.t1.clk  = \AES.r8.t3.clk ;
    assign \AES.r8.t3.t1.in  = \AES.r8.t3.b1 ;
    assign \AES.r8.t3.k1  = \AES.r8.t3.t1.out ;
    assign \AES.r8.t3.t1.s0.clk  = \AES.r8.t3.t1.clk ;
    assign \AES.r8.t3.t1.s0.in  = \AES.r8.t3.t1.in ;
    assign \AES.r8.t3.t1.k0  = \AES.r8.t3.t1.s0.out ;
    always @ (  posedge \AES.r8.t3.t1.s0.clk )
    begin
        case ( \AES.r8.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t1.s4.clk  = \AES.r8.t3.t1.clk ;
    assign \AES.r8.t3.t1.s4.in  = \AES.r8.t3.t1.in ;
    assign \AES.r8.t3.t1.k1  = \AES.r8.t3.t1.s4.out ;
    always @ (  posedge \AES.r8.t3.t1.s4.clk )
    begin
        case ( \AES.r8.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t1.out  = { \AES.r8.t3.t1.k0 , \AES.r8.t3.t1.k0 , ( \AES.r8.t3.t1.k0  ^ \AES.r8.t3.t1.k1  ), \AES.r8.t3.t1.k1  };
    assign \AES.r8.t3.t2.clk  = \AES.r8.t3.clk ;
    assign \AES.r8.t3.t2.in  = \AES.r8.t3.b2 ;
    assign \AES.r8.t3.k2  = \AES.r8.t3.t2.out ;
    assign \AES.r8.t3.t2.s0.clk  = \AES.r8.t3.t2.clk ;
    assign \AES.r8.t3.t2.s0.in  = \AES.r8.t3.t2.in ;
    assign \AES.r8.t3.t2.k0  = \AES.r8.t3.t2.s0.out ;
    always @ (  posedge \AES.r8.t3.t2.s0.clk )
    begin
        case ( \AES.r8.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t2.s4.clk  = \AES.r8.t3.t2.clk ;
    assign \AES.r8.t3.t2.s4.in  = \AES.r8.t3.t2.in ;
    assign \AES.r8.t3.t2.k1  = \AES.r8.t3.t2.s4.out ;
    always @ (  posedge \AES.r8.t3.t2.s4.clk )
    begin
        case ( \AES.r8.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t2.out  = { \AES.r8.t3.t2.k0 , \AES.r8.t3.t2.k0 , ( \AES.r8.t3.t2.k0  ^ \AES.r8.t3.t2.k1  ), \AES.r8.t3.t2.k1  };
    assign \AES.r8.t3.t3.clk  = \AES.r8.t3.clk ;
    assign \AES.r8.t3.t3.in  = \AES.r8.t3.b3 ;
    assign \AES.r8.t3.p3  = \AES.r8.t3.t3.out ;
    assign \AES.r8.t3.t3.s0.clk  = \AES.r8.t3.t3.clk ;
    assign \AES.r8.t3.t3.s0.in  = \AES.r8.t3.t3.in ;
    assign \AES.r8.t3.t3.k0  = \AES.r8.t3.t3.s0.out ;
    always @ (  posedge \AES.r8.t3.t3.s0.clk )
    begin
        case ( \AES.r8.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t3.s4.clk  = \AES.r8.t3.t3.clk ;
    assign \AES.r8.t3.t3.s4.in  = \AES.r8.t3.t3.in ;
    assign \AES.r8.t3.t3.k1  = \AES.r8.t3.t3.s4.out ;
    always @ (  posedge \AES.r8.t3.t3.s4.clk )
    begin
        case ( \AES.r8.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r8.t3.t3.out  = { \AES.r8.t3.t3.k0 , \AES.r8.t3.t3.k0 , ( \AES.r8.t3.t3.k0  ^ \AES.r8.t3.t3.k1  ), \AES.r8.t3.t3.k1  };
    assign \AES.r8.z0  = ( ( ( ( \AES.r8.p00  ^ \AES.r8.p11  ) ^ \AES.r8.p22  ) ^ \AES.r8.p33  ) ^ \AES.r8.k0  );
    assign \AES.r8.z1  = ( ( ( ( \AES.r8.p03  ^ \AES.r8.p10  ) ^ \AES.r8.p21  ) ^ \AES.r8.p32  ) ^ \AES.r8.k1  );
    assign \AES.r8.z2  = ( ( ( ( \AES.r8.p02  ^ \AES.r8.p13  ) ^ \AES.r8.p20  ) ^ \AES.r8.p31  ) ^ \AES.r8.k2  );
    assign \AES.r8.z3  = ( ( ( ( \AES.r8.p01  ^ \AES.r8.p12  ) ^ \AES.r8.p23  ) ^ \AES.r8.p30  ) ^ \AES.r8.k3  );
    always @ (  posedge \AES.r8.clk )
    begin
    end
    assign \AES.r9.clk  = \AES.clk ;
    assign \AES.r9.state_in  = \AES.s8 ;
    assign \AES.r9.key  = \AES.k8b ;
    assign \AES.s9  = \AES.r9.state_out ;
    assign \AES.r9.k0  = \AES.r9.key [127:96];
    assign \AES.r9.k1  = \AES.r9.key [95:64];
    assign \AES.r9.k2  = \AES.r9.key [63:32];
    assign \AES.r9.k3  = \AES.r9.key [31:0];
    assign \AES.r9.s0  = \AES.r9.state_in [127:96];
    assign \AES.r9.s1  = \AES.r9.state_in [95:64];
    assign \AES.r9.s2  = \AES.r9.state_in [63:32];
    assign \AES.r9.s3  = \AES.r9.state_in [31:0];
    assign \AES.r9.t0.clk  = \AES.r9.clk ;
    assign \AES.r9.t0.state  = \AES.r9.s0 ;
    assign \AES.r9.p00  = \AES.r9.t0.p0 ;
    assign \AES.r9.p01  = \AES.r9.t0.p1 ;
    assign \AES.r9.p02  = \AES.r9.t0.p2 ;
    assign \AES.r9.p03  = \AES.r9.t0.p3 ;
    assign \AES.r9.t0.p0  = { \AES.r9.t0.k0 [7:0], \AES.r9.t0.k0 [31:8] };
    assign \AES.r9.t0.p1  = { \AES.r9.t0.k1 [15:0], \AES.r9.t0.k1 [31:16] };
    assign \AES.r9.t0.p2  = { \AES.r9.t0.k2 [23:0], \AES.r9.t0.k2 [31:24] };
    assign \AES.r9.t0.b0  = \AES.r9.t0.state [31:24];
    assign \AES.r9.t0.b1  = \AES.r9.t0.state [23:16];
    assign \AES.r9.t0.b2  = \AES.r9.t0.state [15:8];
    assign \AES.r9.t0.b3  = \AES.r9.t0.state [7:0];
    assign \AES.r9.t0.t0.clk  = \AES.r9.t0.clk ;
    assign \AES.r9.t0.t0.in  = \AES.r9.t0.b0 ;
    assign \AES.r9.t0.k0  = \AES.r9.t0.t0.out ;
    assign \AES.r9.t0.t0.s0.clk  = \AES.r9.t0.t0.clk ;
    assign \AES.r9.t0.t0.s0.in  = \AES.r9.t0.t0.in ;
    assign \AES.r9.t0.t0.k0  = \AES.r9.t0.t0.s0.out ;
    always @ (  posedge \AES.r9.t0.t0.s0.clk )
    begin
        case ( \AES.r9.t0.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t0.s4.clk  = \AES.r9.t0.t0.clk ;
    assign \AES.r9.t0.t0.s4.in  = \AES.r9.t0.t0.in ;
    assign \AES.r9.t0.t0.k1  = \AES.r9.t0.t0.s4.out ;
    always @ (  posedge \AES.r9.t0.t0.s4.clk )
    begin
        case ( \AES.r9.t0.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t0.out  = { \AES.r9.t0.t0.k0 , \AES.r9.t0.t0.k0 , ( \AES.r9.t0.t0.k0  ^ \AES.r9.t0.t0.k1  ), \AES.r9.t0.t0.k1  };
    assign \AES.r9.t0.t1.clk  = \AES.r9.t0.clk ;
    assign \AES.r9.t0.t1.in  = \AES.r9.t0.b1 ;
    assign \AES.r9.t0.k1  = \AES.r9.t0.t1.out ;
    assign \AES.r9.t0.t1.s0.clk  = \AES.r9.t0.t1.clk ;
    assign \AES.r9.t0.t1.s0.in  = \AES.r9.t0.t1.in ;
    assign \AES.r9.t0.t1.k0  = \AES.r9.t0.t1.s0.out ;
    always @ (  posedge \AES.r9.t0.t1.s0.clk )
    begin
        case ( \AES.r9.t0.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t1.s4.clk  = \AES.r9.t0.t1.clk ;
    assign \AES.r9.t0.t1.s4.in  = \AES.r9.t0.t1.in ;
    assign \AES.r9.t0.t1.k1  = \AES.r9.t0.t1.s4.out ;
    always @ (  posedge \AES.r9.t0.t1.s4.clk )
    begin
        case ( \AES.r9.t0.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t1.out  = { \AES.r9.t0.t1.k0 , \AES.r9.t0.t1.k0 , ( \AES.r9.t0.t1.k0  ^ \AES.r9.t0.t1.k1  ), \AES.r9.t0.t1.k1  };
    assign \AES.r9.t0.t2.clk  = \AES.r9.t0.clk ;
    assign \AES.r9.t0.t2.in  = \AES.r9.t0.b2 ;
    assign \AES.r9.t0.k2  = \AES.r9.t0.t2.out ;
    assign \AES.r9.t0.t2.s0.clk  = \AES.r9.t0.t2.clk ;
    assign \AES.r9.t0.t2.s0.in  = \AES.r9.t0.t2.in ;
    assign \AES.r9.t0.t2.k0  = \AES.r9.t0.t2.s0.out ;
    always @ (  posedge \AES.r9.t0.t2.s0.clk )
    begin
        case ( \AES.r9.t0.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t2.s4.clk  = \AES.r9.t0.t2.clk ;
    assign \AES.r9.t0.t2.s4.in  = \AES.r9.t0.t2.in ;
    assign \AES.r9.t0.t2.k1  = \AES.r9.t0.t2.s4.out ;
    always @ (  posedge \AES.r9.t0.t2.s4.clk )
    begin
        case ( \AES.r9.t0.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t2.out  = { \AES.r9.t0.t2.k0 , \AES.r9.t0.t2.k0 , ( \AES.r9.t0.t2.k0  ^ \AES.r9.t0.t2.k1  ), \AES.r9.t0.t2.k1  };
    assign \AES.r9.t0.t3.clk  = \AES.r9.t0.clk ;
    assign \AES.r9.t0.t3.in  = \AES.r9.t0.b3 ;
    assign \AES.r9.t0.p3  = \AES.r9.t0.t3.out ;
    assign \AES.r9.t0.t3.s0.clk  = \AES.r9.t0.t3.clk ;
    assign \AES.r9.t0.t3.s0.in  = \AES.r9.t0.t3.in ;
    assign \AES.r9.t0.t3.k0  = \AES.r9.t0.t3.s0.out ;
    always @ (  posedge \AES.r9.t0.t3.s0.clk )
    begin
        case ( \AES.r9.t0.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t3.s4.clk  = \AES.r9.t0.t3.clk ;
    assign \AES.r9.t0.t3.s4.in  = \AES.r9.t0.t3.in ;
    assign \AES.r9.t0.t3.k1  = \AES.r9.t0.t3.s4.out ;
    always @ (  posedge \AES.r9.t0.t3.s4.clk )
    begin
        case ( \AES.r9.t0.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t0.t3.out  = { \AES.r9.t0.t3.k0 , \AES.r9.t0.t3.k0 , ( \AES.r9.t0.t3.k0  ^ \AES.r9.t0.t3.k1  ), \AES.r9.t0.t3.k1  };
    assign \AES.r9.t1.clk  = \AES.r9.clk ;
    assign \AES.r9.t1.state  = \AES.r9.s1 ;
    assign \AES.r9.p10  = \AES.r9.t1.p0 ;
    assign \AES.r9.p11  = \AES.r9.t1.p1 ;
    assign \AES.r9.p12  = \AES.r9.t1.p2 ;
    assign \AES.r9.p13  = \AES.r9.t1.p3 ;
    assign \AES.r9.t1.p0  = { \AES.r9.t1.k0 [7:0], \AES.r9.t1.k0 [31:8] };
    assign \AES.r9.t1.p1  = { \AES.r9.t1.k1 [15:0], \AES.r9.t1.k1 [31:16] };
    assign \AES.r9.t1.p2  = { \AES.r9.t1.k2 [23:0], \AES.r9.t1.k2 [31:24] };
    assign \AES.r9.t1.b0  = \AES.r9.t1.state [31:24];
    assign \AES.r9.t1.b1  = \AES.r9.t1.state [23:16];
    assign \AES.r9.t1.b2  = \AES.r9.t1.state [15:8];
    assign \AES.r9.t1.b3  = \AES.r9.t1.state [7:0];
    assign \AES.r9.t1.t0.clk  = \AES.r9.t1.clk ;
    assign \AES.r9.t1.t0.in  = \AES.r9.t1.b0 ;
    assign \AES.r9.t1.k0  = \AES.r9.t1.t0.out ;
    assign \AES.r9.t1.t0.s0.clk  = \AES.r9.t1.t0.clk ;
    assign \AES.r9.t1.t0.s0.in  = \AES.r9.t1.t0.in ;
    assign \AES.r9.t1.t0.k0  = \AES.r9.t1.t0.s0.out ;
    always @ (  posedge \AES.r9.t1.t0.s0.clk )
    begin
        case ( \AES.r9.t1.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t0.s4.clk  = \AES.r9.t1.t0.clk ;
    assign \AES.r9.t1.t0.s4.in  = \AES.r9.t1.t0.in ;
    assign \AES.r9.t1.t0.k1  = \AES.r9.t1.t0.s4.out ;
    always @ (  posedge \AES.r9.t1.t0.s4.clk )
    begin
        case ( \AES.r9.t1.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t0.out  = { \AES.r9.t1.t0.k0 , \AES.r9.t1.t0.k0 , ( \AES.r9.t1.t0.k0  ^ \AES.r9.t1.t0.k1  ), \AES.r9.t1.t0.k1  };
    assign \AES.r9.t1.t1.clk  = \AES.r9.t1.clk ;
    assign \AES.r9.t1.t1.in  = \AES.r9.t1.b1 ;
    assign \AES.r9.t1.k1  = \AES.r9.t1.t1.out ;
    assign \AES.r9.t1.t1.s0.clk  = \AES.r9.t1.t1.clk ;
    assign \AES.r9.t1.t1.s0.in  = \AES.r9.t1.t1.in ;
    assign \AES.r9.t1.t1.k0  = \AES.r9.t1.t1.s0.out ;
    always @ (  posedge \AES.r9.t1.t1.s0.clk )
    begin
        case ( \AES.r9.t1.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t1.s4.clk  = \AES.r9.t1.t1.clk ;
    assign \AES.r9.t1.t1.s4.in  = \AES.r9.t1.t1.in ;
    assign \AES.r9.t1.t1.k1  = \AES.r9.t1.t1.s4.out ;
    always @ (  posedge \AES.r9.t1.t1.s4.clk )
    begin
        case ( \AES.r9.t1.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t1.out  = { \AES.r9.t1.t1.k0 , \AES.r9.t1.t1.k0 , ( \AES.r9.t1.t1.k0  ^ \AES.r9.t1.t1.k1  ), \AES.r9.t1.t1.k1  };
    assign \AES.r9.t1.t2.clk  = \AES.r9.t1.clk ;
    assign \AES.r9.t1.t2.in  = \AES.r9.t1.b2 ;
    assign \AES.r9.t1.k2  = \AES.r9.t1.t2.out ;
    assign \AES.r9.t1.t2.s0.clk  = \AES.r9.t1.t2.clk ;
    assign \AES.r9.t1.t2.s0.in  = \AES.r9.t1.t2.in ;
    assign \AES.r9.t1.t2.k0  = \AES.r9.t1.t2.s0.out ;
    always @ (  posedge \AES.r9.t1.t2.s0.clk )
    begin
        case ( \AES.r9.t1.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t2.s4.clk  = \AES.r9.t1.t2.clk ;
    assign \AES.r9.t1.t2.s4.in  = \AES.r9.t1.t2.in ;
    assign \AES.r9.t1.t2.k1  = \AES.r9.t1.t2.s4.out ;
    always @ (  posedge \AES.r9.t1.t2.s4.clk )
    begin
        case ( \AES.r9.t1.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t2.out  = { \AES.r9.t1.t2.k0 , \AES.r9.t1.t2.k0 , ( \AES.r9.t1.t2.k0  ^ \AES.r9.t1.t2.k1  ), \AES.r9.t1.t2.k1  };
    assign \AES.r9.t1.t3.clk  = \AES.r9.t1.clk ;
    assign \AES.r9.t1.t3.in  = \AES.r9.t1.b3 ;
    assign \AES.r9.t1.p3  = \AES.r9.t1.t3.out ;
    assign \AES.r9.t1.t3.s0.clk  = \AES.r9.t1.t3.clk ;
    assign \AES.r9.t1.t3.s0.in  = \AES.r9.t1.t3.in ;
    assign \AES.r9.t1.t3.k0  = \AES.r9.t1.t3.s0.out ;
    always @ (  posedge \AES.r9.t1.t3.s0.clk )
    begin
        case ( \AES.r9.t1.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t3.s4.clk  = \AES.r9.t1.t3.clk ;
    assign \AES.r9.t1.t3.s4.in  = \AES.r9.t1.t3.in ;
    assign \AES.r9.t1.t3.k1  = \AES.r9.t1.t3.s4.out ;
    always @ (  posedge \AES.r9.t1.t3.s4.clk )
    begin
        case ( \AES.r9.t1.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t1.t3.out  = { \AES.r9.t1.t3.k0 , \AES.r9.t1.t3.k0 , ( \AES.r9.t1.t3.k0  ^ \AES.r9.t1.t3.k1  ), \AES.r9.t1.t3.k1  };
    assign \AES.r9.t2.clk  = \AES.r9.clk ;
    assign \AES.r9.t2.state  = \AES.r9.s2 ;
    assign \AES.r9.p20  = \AES.r9.t2.p0 ;
    assign \AES.r9.p21  = \AES.r9.t2.p1 ;
    assign \AES.r9.p22  = \AES.r9.t2.p2 ;
    assign \AES.r9.p23  = \AES.r9.t2.p3 ;
    assign \AES.r9.t2.p0  = { \AES.r9.t2.k0 [7:0], \AES.r9.t2.k0 [31:8] };
    assign \AES.r9.t2.p1  = { \AES.r9.t2.k1 [15:0], \AES.r9.t2.k1 [31:16] };
    assign \AES.r9.t2.p2  = { \AES.r9.t2.k2 [23:0], \AES.r9.t2.k2 [31:24] };
    assign \AES.r9.t2.b0  = \AES.r9.t2.state [31:24];
    assign \AES.r9.t2.b1  = \AES.r9.t2.state [23:16];
    assign \AES.r9.t2.b2  = \AES.r9.t2.state [15:8];
    assign \AES.r9.t2.b3  = \AES.r9.t2.state [7:0];
    assign \AES.r9.t2.t0.clk  = \AES.r9.t2.clk ;
    assign \AES.r9.t2.t0.in  = \AES.r9.t2.b0 ;
    assign \AES.r9.t2.k0  = \AES.r9.t2.t0.out ;
    assign \AES.r9.t2.t0.s0.clk  = \AES.r9.t2.t0.clk ;
    assign \AES.r9.t2.t0.s0.in  = \AES.r9.t2.t0.in ;
    assign \AES.r9.t2.t0.k0  = \AES.r9.t2.t0.s0.out ;
    always @ (  posedge \AES.r9.t2.t0.s0.clk )
    begin
        case ( \AES.r9.t2.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t0.s4.clk  = \AES.r9.t2.t0.clk ;
    assign \AES.r9.t2.t0.s4.in  = \AES.r9.t2.t0.in ;
    assign \AES.r9.t2.t0.k1  = \AES.r9.t2.t0.s4.out ;
    always @ (  posedge \AES.r9.t2.t0.s4.clk )
    begin
        case ( \AES.r9.t2.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t0.out  = { \AES.r9.t2.t0.k0 , \AES.r9.t2.t0.k0 , ( \AES.r9.t2.t0.k0  ^ \AES.r9.t2.t0.k1  ), \AES.r9.t2.t0.k1  };
    assign \AES.r9.t2.t1.clk  = \AES.r9.t2.clk ;
    assign \AES.r9.t2.t1.in  = \AES.r9.t2.b1 ;
    assign \AES.r9.t2.k1  = \AES.r9.t2.t1.out ;
    assign \AES.r9.t2.t1.s0.clk  = \AES.r9.t2.t1.clk ;
    assign \AES.r9.t2.t1.s0.in  = \AES.r9.t2.t1.in ;
    assign \AES.r9.t2.t1.k0  = \AES.r9.t2.t1.s0.out ;
    always @ (  posedge \AES.r9.t2.t1.s0.clk )
    begin
        case ( \AES.r9.t2.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t1.s4.clk  = \AES.r9.t2.t1.clk ;
    assign \AES.r9.t2.t1.s4.in  = \AES.r9.t2.t1.in ;
    assign \AES.r9.t2.t1.k1  = \AES.r9.t2.t1.s4.out ;
    always @ (  posedge \AES.r9.t2.t1.s4.clk )
    begin
        case ( \AES.r9.t2.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t1.out  = { \AES.r9.t2.t1.k0 , \AES.r9.t2.t1.k0 , ( \AES.r9.t2.t1.k0  ^ \AES.r9.t2.t1.k1  ), \AES.r9.t2.t1.k1  };
    assign \AES.r9.t2.t2.clk  = \AES.r9.t2.clk ;
    assign \AES.r9.t2.t2.in  = \AES.r9.t2.b2 ;
    assign \AES.r9.t2.k2  = \AES.r9.t2.t2.out ;
    assign \AES.r9.t2.t2.s0.clk  = \AES.r9.t2.t2.clk ;
    assign \AES.r9.t2.t2.s0.in  = \AES.r9.t2.t2.in ;
    assign \AES.r9.t2.t2.k0  = \AES.r9.t2.t2.s0.out ;
    always @ (  posedge \AES.r9.t2.t2.s0.clk )
    begin
        case ( \AES.r9.t2.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t2.s4.clk  = \AES.r9.t2.t2.clk ;
    assign \AES.r9.t2.t2.s4.in  = \AES.r9.t2.t2.in ;
    assign \AES.r9.t2.t2.k1  = \AES.r9.t2.t2.s4.out ;
    always @ (  posedge \AES.r9.t2.t2.s4.clk )
    begin
        case ( \AES.r9.t2.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t2.out  = { \AES.r9.t2.t2.k0 , \AES.r9.t2.t2.k0 , ( \AES.r9.t2.t2.k0  ^ \AES.r9.t2.t2.k1  ), \AES.r9.t2.t2.k1  };
    assign \AES.r9.t2.t3.clk  = \AES.r9.t2.clk ;
    assign \AES.r9.t2.t3.in  = \AES.r9.t2.b3 ;
    assign \AES.r9.t2.p3  = \AES.r9.t2.t3.out ;
    assign \AES.r9.t2.t3.s0.clk  = \AES.r9.t2.t3.clk ;
    assign \AES.r9.t2.t3.s0.in  = \AES.r9.t2.t3.in ;
    assign \AES.r9.t2.t3.k0  = \AES.r9.t2.t3.s0.out ;
    always @ (  posedge \AES.r9.t2.t3.s0.clk )
    begin
        case ( \AES.r9.t2.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t3.s4.clk  = \AES.r9.t2.t3.clk ;
    assign \AES.r9.t2.t3.s4.in  = \AES.r9.t2.t3.in ;
    assign \AES.r9.t2.t3.k1  = \AES.r9.t2.t3.s4.out ;
    always @ (  posedge \AES.r9.t2.t3.s4.clk )
    begin
        case ( \AES.r9.t2.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t2.t3.out  = { \AES.r9.t2.t3.k0 , \AES.r9.t2.t3.k0 , ( \AES.r9.t2.t3.k0  ^ \AES.r9.t2.t3.k1  ), \AES.r9.t2.t3.k1  };
    assign \AES.r9.t3.clk  = \AES.r9.clk ;
    assign \AES.r9.t3.state  = \AES.r9.s3 ;
    assign \AES.r9.p30  = \AES.r9.t3.p0 ;
    assign \AES.r9.p31  = \AES.r9.t3.p1 ;
    assign \AES.r9.p32  = \AES.r9.t3.p2 ;
    assign \AES.r9.p33  = \AES.r9.t3.p3 ;
    assign \AES.r9.t3.p0  = { \AES.r9.t3.k0 [7:0], \AES.r9.t3.k0 [31:8] };
    assign \AES.r9.t3.p1  = { \AES.r9.t3.k1 [15:0], \AES.r9.t3.k1 [31:16] };
    assign \AES.r9.t3.p2  = { \AES.r9.t3.k2 [23:0], \AES.r9.t3.k2 [31:24] };
    assign \AES.r9.t3.b0  = \AES.r9.t3.state [31:24];
    assign \AES.r9.t3.b1  = \AES.r9.t3.state [23:16];
    assign \AES.r9.t3.b2  = \AES.r9.t3.state [15:8];
    assign \AES.r9.t3.b3  = \AES.r9.t3.state [7:0];
    assign \AES.r9.t3.t0.clk  = \AES.r9.t3.clk ;
    assign \AES.r9.t3.t0.in  = \AES.r9.t3.b0 ;
    assign \AES.r9.t3.k0  = \AES.r9.t3.t0.out ;
    assign \AES.r9.t3.t0.s0.clk  = \AES.r9.t3.t0.clk ;
    assign \AES.r9.t3.t0.s0.in  = \AES.r9.t3.t0.in ;
    assign \AES.r9.t3.t0.k0  = \AES.r9.t3.t0.s0.out ;
    always @ (  posedge \AES.r9.t3.t0.s0.clk )
    begin
        case ( \AES.r9.t3.t0.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t0.s4.clk  = \AES.r9.t3.t0.clk ;
    assign \AES.r9.t3.t0.s4.in  = \AES.r9.t3.t0.in ;
    assign \AES.r9.t3.t0.k1  = \AES.r9.t3.t0.s4.out ;
    always @ (  posedge \AES.r9.t3.t0.s4.clk )
    begin
        case ( \AES.r9.t3.t0.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t0.out  = { \AES.r9.t3.t0.k0 , \AES.r9.t3.t0.k0 , ( \AES.r9.t3.t0.k0  ^ \AES.r9.t3.t0.k1  ), \AES.r9.t3.t0.k1  };
    assign \AES.r9.t3.t1.clk  = \AES.r9.t3.clk ;
    assign \AES.r9.t3.t1.in  = \AES.r9.t3.b1 ;
    assign \AES.r9.t3.k1  = \AES.r9.t3.t1.out ;
    assign \AES.r9.t3.t1.s0.clk  = \AES.r9.t3.t1.clk ;
    assign \AES.r9.t3.t1.s0.in  = \AES.r9.t3.t1.in ;
    assign \AES.r9.t3.t1.k0  = \AES.r9.t3.t1.s0.out ;
    always @ (  posedge \AES.r9.t3.t1.s0.clk )
    begin
        case ( \AES.r9.t3.t1.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t1.s4.clk  = \AES.r9.t3.t1.clk ;
    assign \AES.r9.t3.t1.s4.in  = \AES.r9.t3.t1.in ;
    assign \AES.r9.t3.t1.k1  = \AES.r9.t3.t1.s4.out ;
    always @ (  posedge \AES.r9.t3.t1.s4.clk )
    begin
        case ( \AES.r9.t3.t1.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t1.out  = { \AES.r9.t3.t1.k0 , \AES.r9.t3.t1.k0 , ( \AES.r9.t3.t1.k0  ^ \AES.r9.t3.t1.k1  ), \AES.r9.t3.t1.k1  };
    assign \AES.r9.t3.t2.clk  = \AES.r9.t3.clk ;
    assign \AES.r9.t3.t2.in  = \AES.r9.t3.b2 ;
    assign \AES.r9.t3.k2  = \AES.r9.t3.t2.out ;
    assign \AES.r9.t3.t2.s0.clk  = \AES.r9.t3.t2.clk ;
    assign \AES.r9.t3.t2.s0.in  = \AES.r9.t3.t2.in ;
    assign \AES.r9.t3.t2.k0  = \AES.r9.t3.t2.s0.out ;
    always @ (  posedge \AES.r9.t3.t2.s0.clk )
    begin
        case ( \AES.r9.t3.t2.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t2.s4.clk  = \AES.r9.t3.t2.clk ;
    assign \AES.r9.t3.t2.s4.in  = \AES.r9.t3.t2.in ;
    assign \AES.r9.t3.t2.k1  = \AES.r9.t3.t2.s4.out ;
    always @ (  posedge \AES.r9.t3.t2.s4.clk )
    begin
        case ( \AES.r9.t3.t2.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t2.out  = { \AES.r9.t3.t2.k0 , \AES.r9.t3.t2.k0 , ( \AES.r9.t3.t2.k0  ^ \AES.r9.t3.t2.k1  ), \AES.r9.t3.t2.k1  };
    assign \AES.r9.t3.t3.clk  = \AES.r9.t3.clk ;
    assign \AES.r9.t3.t3.in  = \AES.r9.t3.b3 ;
    assign \AES.r9.t3.p3  = \AES.r9.t3.t3.out ;
    assign \AES.r9.t3.t3.s0.clk  = \AES.r9.t3.t3.clk ;
    assign \AES.r9.t3.t3.s0.in  = \AES.r9.t3.t3.in ;
    assign \AES.r9.t3.t3.k0  = \AES.r9.t3.t3.s0.out ;
    always @ (  posedge \AES.r9.t3.t3.s0.clk )
    begin
        case ( \AES.r9.t3.t3.s0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t3.s4.clk  = \AES.r9.t3.t3.clk ;
    assign \AES.r9.t3.t3.s4.in  = \AES.r9.t3.t3.in ;
    assign \AES.r9.t3.t3.k1  = \AES.r9.t3.t3.s4.out ;
    always @ (  posedge \AES.r9.t3.t3.s4.clk )
    begin
        case ( \AES.r9.t3.t3.s4.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.r9.t3.t3.out  = { \AES.r9.t3.t3.k0 , \AES.r9.t3.t3.k0 , ( \AES.r9.t3.t3.k0  ^ \AES.r9.t3.t3.k1  ), \AES.r9.t3.t3.k1  };
    assign \AES.r9.z0  = ( ( ( ( \AES.r9.p00  ^ \AES.r9.p11  ) ^ \AES.r9.p22  ) ^ \AES.r9.p33  ) ^ \AES.r9.k0  );
    assign \AES.r9.z1  = ( ( ( ( \AES.r9.p03  ^ \AES.r9.p10  ) ^ \AES.r9.p21  ) ^ \AES.r9.p32  ) ^ \AES.r9.k1  );
    assign \AES.r9.z2  = ( ( ( ( \AES.r9.p02  ^ \AES.r9.p13  ) ^ \AES.r9.p20  ) ^ \AES.r9.p31  ) ^ \AES.r9.k2  );
    assign \AES.r9.z3  = ( ( ( ( \AES.r9.p01  ^ \AES.r9.p12  ) ^ \AES.r9.p23  ) ^ \AES.r9.p30  ) ^ \AES.r9.k3  );
    always @ (  posedge \AES.r9.clk )
    begin
    end
    assign \AES.rf.clk  = \AES.clk ;
    assign \AES.rf.state_in  = \AES.s9 ;
    assign \AES.rf.key_in  = \AES.k9b ;
    assign \AES.out  = \AES.rf.state_out ;
    assign \AES.rf.k0  = \AES.rf.key_in [127:96];
    assign \AES.rf.k1  = \AES.rf.key_in [95:64];
    assign \AES.rf.k2  = \AES.rf.key_in [63:32];
    assign \AES.rf.k3  = \AES.rf.key_in [31:0];
    assign \AES.rf.s0  = \AES.rf.state_in [127:96];
    assign \AES.rf.s1  = \AES.rf.state_in [95:64];
    assign \AES.rf.s2  = \AES.rf.state_in [63:32];
    assign \AES.rf.s3  = \AES.rf.state_in [31:0];
    assign \AES.rf.S4_1.clk  = \AES.rf.clk ;
    assign \AES.rf.S4_1.in  = \AES.rf.s0 ;
    assign \AES.rf.S4_1.S_0.clk  = \AES.rf.S4_1.clk ;
    assign \AES.rf.S4_1.S_0.in  = \AES.rf.S4_1.in [31:24];
    assign \AES.rf.S4_1.k0  = \AES.rf.S4_1.S_0.out ;
    always @ (  posedge \AES.rf.S4_1.S_0.clk )
    begin
        case ( \AES.rf.S4_1.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_1.S_1.clk  = \AES.rf.S4_1.clk ;
    assign \AES.rf.S4_1.S_1.in  = \AES.rf.S4_1.in [23:16];
    assign \AES.rf.S4_1.k1  = \AES.rf.S4_1.S_1.out ;
    always @ (  posedge \AES.rf.S4_1.S_1.clk )
    begin
        case ( \AES.rf.S4_1.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_1.S_2.clk  = \AES.rf.S4_1.clk ;
    assign \AES.rf.S4_1.S_2.in  = \AES.rf.S4_1.in [15:8];
    assign \AES.rf.S4_1.k2  = \AES.rf.S4_1.S_2.out ;
    always @ (  posedge \AES.rf.S4_1.S_2.clk )
    begin
        case ( \AES.rf.S4_1.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_1.S_3.clk  = \AES.rf.S4_1.clk ;
    assign \AES.rf.S4_1.S_3.in  = \AES.rf.S4_1.in [7:0];
    assign \AES.rf.S4_1.k3  = \AES.rf.S4_1.S_3.out ;
    always @ (  posedge \AES.rf.S4_1.S_3.clk )
    begin
        case ( \AES.rf.S4_1.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_1.out  = { \AES.rf.S4_1.k0 , \AES.rf.S4_1.k1 , \AES.rf.S4_1.k2 , \AES.rf.S4_1.k3  };
    assign \AES.rf.S4_2.clk  = \AES.rf.clk ;
    assign \AES.rf.S4_2.in  = \AES.rf.s1 ;
    assign \AES.rf.S4_2.S_0.clk  = \AES.rf.S4_2.clk ;
    assign \AES.rf.S4_2.S_0.in  = \AES.rf.S4_2.in [31:24];
    assign \AES.rf.S4_2.k0  = \AES.rf.S4_2.S_0.out ;
    always @ (  posedge \AES.rf.S4_2.S_0.clk )
    begin
        case ( \AES.rf.S4_2.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_2.S_1.clk  = \AES.rf.S4_2.clk ;
    assign \AES.rf.S4_2.S_1.in  = \AES.rf.S4_2.in [23:16];
    assign \AES.rf.S4_2.k1  = \AES.rf.S4_2.S_1.out ;
    always @ (  posedge \AES.rf.S4_2.S_1.clk )
    begin
        case ( \AES.rf.S4_2.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_2.S_2.clk  = \AES.rf.S4_2.clk ;
    assign \AES.rf.S4_2.S_2.in  = \AES.rf.S4_2.in [15:8];
    assign \AES.rf.S4_2.k2  = \AES.rf.S4_2.S_2.out ;
    always @ (  posedge \AES.rf.S4_2.S_2.clk )
    begin
        case ( \AES.rf.S4_2.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_2.S_3.clk  = \AES.rf.S4_2.clk ;
    assign \AES.rf.S4_2.S_3.in  = \AES.rf.S4_2.in [7:0];
    assign \AES.rf.S4_2.k3  = \AES.rf.S4_2.S_3.out ;
    always @ (  posedge \AES.rf.S4_2.S_3.clk )
    begin
        case ( \AES.rf.S4_2.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_2.out  = { \AES.rf.S4_2.k0 , \AES.rf.S4_2.k1 , \AES.rf.S4_2.k2 , \AES.rf.S4_2.k3  };
    assign \AES.rf.S4_3.clk  = \AES.rf.clk ;
    assign \AES.rf.S4_3.in  = \AES.rf.s2 ;
    assign \AES.rf.S4_3.S_0.clk  = \AES.rf.S4_3.clk ;
    assign \AES.rf.S4_3.S_0.in  = \AES.rf.S4_3.in [31:24];
    assign \AES.rf.S4_3.k0  = \AES.rf.S4_3.S_0.out ;
    always @ (  posedge \AES.rf.S4_3.S_0.clk )
    begin
        case ( \AES.rf.S4_3.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_3.S_1.clk  = \AES.rf.S4_3.clk ;
    assign \AES.rf.S4_3.S_1.in  = \AES.rf.S4_3.in [23:16];
    assign \AES.rf.S4_3.k1  = \AES.rf.S4_3.S_1.out ;
    always @ (  posedge \AES.rf.S4_3.S_1.clk )
    begin
        case ( \AES.rf.S4_3.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_3.S_2.clk  = \AES.rf.S4_3.clk ;
    assign \AES.rf.S4_3.S_2.in  = \AES.rf.S4_3.in [15:8];
    assign \AES.rf.S4_3.k2  = \AES.rf.S4_3.S_2.out ;
    always @ (  posedge \AES.rf.S4_3.S_2.clk )
    begin
        case ( \AES.rf.S4_3.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_3.S_3.clk  = \AES.rf.S4_3.clk ;
    assign \AES.rf.S4_3.S_3.in  = \AES.rf.S4_3.in [7:0];
    assign \AES.rf.S4_3.k3  = \AES.rf.S4_3.S_3.out ;
    always @ (  posedge \AES.rf.S4_3.S_3.clk )
    begin
        case ( \AES.rf.S4_3.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_3.out  = { \AES.rf.S4_3.k0 , \AES.rf.S4_3.k1 , \AES.rf.S4_3.k2 , \AES.rf.S4_3.k3  };
    assign \AES.rf.S4_4.clk  = \AES.rf.clk ;
    assign \AES.rf.S4_4.in  = \AES.rf.s3 ;
    assign \AES.rf.S4_4.S_0.clk  = \AES.rf.S4_4.clk ;
    assign \AES.rf.S4_4.S_0.in  = \AES.rf.S4_4.in [31:24];
    assign \AES.rf.S4_4.k0  = \AES.rf.S4_4.S_0.out ;
    always @ (  posedge \AES.rf.S4_4.S_0.clk )
    begin
        case ( \AES.rf.S4_4.S_0.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_4.S_1.clk  = \AES.rf.S4_4.clk ;
    assign \AES.rf.S4_4.S_1.in  = \AES.rf.S4_4.in [23:16];
    assign \AES.rf.S4_4.k1  = \AES.rf.S4_4.S_1.out ;
    always @ (  posedge \AES.rf.S4_4.S_1.clk )
    begin
        case ( \AES.rf.S4_4.S_1.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_4.S_2.clk  = \AES.rf.S4_4.clk ;
    assign \AES.rf.S4_4.S_2.in  = \AES.rf.S4_4.in [15:8];
    assign \AES.rf.S4_4.k2  = \AES.rf.S4_4.S_2.out ;
    always @ (  posedge \AES.rf.S4_4.S_2.clk )
    begin
        case ( \AES.rf.S4_4.S_2.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_4.S_3.clk  = \AES.rf.S4_4.clk ;
    assign \AES.rf.S4_4.S_3.in  = \AES.rf.S4_4.in [7:0];
    assign \AES.rf.S4_4.k3  = \AES.rf.S4_4.S_3.out ;
    always @ (  posedge \AES.rf.S4_4.S_3.clk )
    begin
        case ( \AES.rf.S4_4.S_3.in  ) 
        8'h00:
        begin
        end
        8'h01:
        begin
        end
        8'h02:
        begin
        end
        8'h03:
        begin
        end
        8'h04:
        begin
        end
        8'h05:
        begin
        end
        8'h06:
        begin
        end
        8'h07:
        begin
        end
        8'h08:
        begin
        end
        8'h09:
        begin
        end
        8'h0a:
        begin
        end
        8'h0b:
        begin
        end
        8'h0c:
        begin
        end
        8'h0d:
        begin
        end
        8'h0e:
        begin
        end
        8'h0f:
        begin
        end
        8'h10:
        begin
        end
        8'h11:
        begin
        end
        8'h12:
        begin
        end
        8'h13:
        begin
        end
        8'h14:
        begin
        end
        8'h15:
        begin
        end
        8'h16:
        begin
        end
        8'h17:
        begin
        end
        8'h18:
        begin
        end
        8'h19:
        begin
        end
        8'h1a:
        begin
        end
        8'h1b:
        begin
        end
        8'h1c:
        begin
        end
        8'h1d:
        begin
        end
        8'h1e:
        begin
        end
        8'h1f:
        begin
        end
        8'h20:
        begin
        end
        8'h21:
        begin
        end
        8'h22:
        begin
        end
        8'h23:
        begin
        end
        8'h24:
        begin
        end
        8'h25:
        begin
        end
        8'h26:
        begin
        end
        8'h27:
        begin
        end
        8'h28:
        begin
        end
        8'h29:
        begin
        end
        8'h2a:
        begin
        end
        8'h2b:
        begin
        end
        8'h2c:
        begin
        end
        8'h2d:
        begin
        end
        8'h2e:
        begin
        end
        8'h2f:
        begin
        end
        8'h30:
        begin
        end
        8'h31:
        begin
        end
        8'h32:
        begin
        end
        8'h33:
        begin
        end
        8'h34:
        begin
        end
        8'h35:
        begin
        end
        8'h36:
        begin
        end
        8'h37:
        begin
        end
        8'h38:
        begin
        end
        8'h39:
        begin
        end
        8'h3a:
        begin
        end
        8'h3b:
        begin
        end
        8'h3c:
        begin
        end
        8'h3d:
        begin
        end
        8'h3e:
        begin
        end
        8'h3f:
        begin
        end
        8'h40:
        begin
        end
        8'h41:
        begin
        end
        8'h42:
        begin
        end
        8'h43:
        begin
        end
        8'h44:
        begin
        end
        8'h45:
        begin
        end
        8'h46:
        begin
        end
        8'h47:
        begin
        end
        8'h48:
        begin
        end
        8'h49:
        begin
        end
        8'h4a:
        begin
        end
        8'h4b:
        begin
        end
        8'h4c:
        begin
        end
        8'h4d:
        begin
        end
        8'h4e:
        begin
        end
        8'h4f:
        begin
        end
        8'h50:
        begin
        end
        8'h51:
        begin
        end
        8'h52:
        begin
        end
        8'h53:
        begin
        end
        8'h54:
        begin
        end
        8'h55:
        begin
        end
        8'h56:
        begin
        end
        8'h57:
        begin
        end
        8'h58:
        begin
        end
        8'h59:
        begin
        end
        8'h5a:
        begin
        end
        8'h5b:
        begin
        end
        8'h5c:
        begin
        end
        8'h5d:
        begin
        end
        8'h5e:
        begin
        end
        8'h5f:
        begin
        end
        8'h60:
        begin
        end
        8'h61:
        begin
        end
        8'h62:
        begin
        end
        8'h63:
        begin
        end
        8'h64:
        begin
        end
        8'h65:
        begin
        end
        8'h66:
        begin
        end
        8'h67:
        begin
        end
        8'h68:
        begin
        end
        8'h69:
        begin
        end
        8'h6a:
        begin
        end
        8'h6b:
        begin
        end
        8'h6c:
        begin
        end
        8'h6d:
        begin
        end
        8'h6e:
        begin
        end
        8'h6f:
        begin
        end
        8'h70:
        begin
        end
        8'h71:
        begin
        end
        8'h72:
        begin
        end
        8'h73:
        begin
        end
        8'h74:
        begin
        end
        8'h75:
        begin
        end
        8'h76:
        begin
        end
        8'h77:
        begin
        end
        8'h78:
        begin
        end
        8'h79:
        begin
        end
        8'h7a:
        begin
        end
        8'h7b:
        begin
        end
        8'h7c:
        begin
        end
        8'h7d:
        begin
        end
        8'h7e:
        begin
        end
        8'h7f:
        begin
        end
        8'h80:
        begin
        end
        8'h81:
        begin
        end
        8'h82:
        begin
        end
        8'h83:
        begin
        end
        8'h84:
        begin
        end
        8'h85:
        begin
        end
        8'h86:
        begin
        end
        8'h87:
        begin
        end
        8'h88:
        begin
        end
        8'h89:
        begin
        end
        8'h8a:
        begin
        end
        8'h8b:
        begin
        end
        8'h8c:
        begin
        end
        8'h8d:
        begin
        end
        8'h8e:
        begin
        end
        8'h8f:
        begin
        end
        8'h90:
        begin
        end
        8'h91:
        begin
        end
        8'h92:
        begin
        end
        8'h93:
        begin
        end
        8'h94:
        begin
        end
        8'h95:
        begin
        end
        8'h96:
        begin
        end
        8'h97:
        begin
        end
        8'h98:
        begin
        end
        8'h99:
        begin
        end
        8'h9a:
        begin
        end
        8'h9b:
        begin
        end
        8'h9c:
        begin
        end
        8'h9d:
        begin
        end
        8'h9e:
        begin
        end
        8'h9f:
        begin
        end
        8'ha0:
        begin
        end
        8'ha1:
        begin
        end
        8'ha2:
        begin
        end
        8'ha3:
        begin
        end
        8'ha4:
        begin
        end
        8'ha5:
        begin
        end
        8'ha6:
        begin
        end
        8'ha7:
        begin
        end
        8'ha8:
        begin
        end
        8'ha9:
        begin
        end
        8'haa:
        begin
        end
        8'hab:
        begin
        end
        8'hac:
        begin
        end
        8'had:
        begin
        end
        8'hae:
        begin
        end
        8'haf:
        begin
        end
        8'hb0:
        begin
        end
        8'hb1:
        begin
        end
        8'hb2:
        begin
        end
        8'hb3:
        begin
        end
        8'hb4:
        begin
        end
        8'hb5:
        begin
        end
        8'hb6:
        begin
        end
        8'hb7:
        begin
        end
        8'hb8:
        begin
        end
        8'hb9:
        begin
        end
        8'hba:
        begin
        end
        8'hbb:
        begin
        end
        8'hbc:
        begin
        end
        8'hbd:
        begin
        end
        8'hbe:
        begin
        end
        8'hbf:
        begin
        end
        8'hc0:
        begin
        end
        8'hc1:
        begin
        end
        8'hc2:
        begin
        end
        8'hc3:
        begin
        end
        8'hc4:
        begin
        end
        8'hc5:
        begin
        end
        8'hc6:
        begin
        end
        8'hc7:
        begin
        end
        8'hc8:
        begin
        end
        8'hc9:
        begin
        end
        8'hca:
        begin
        end
        8'hcb:
        begin
        end
        8'hcc:
        begin
        end
        8'hcd:
        begin
        end
        8'hce:
        begin
        end
        8'hcf:
        begin
        end
        8'hd0:
        begin
        end
        8'hd1:
        begin
        end
        8'hd2:
        begin
        end
        8'hd3:
        begin
        end
        8'hd4:
        begin
        end
        8'hd5:
        begin
        end
        8'hd6:
        begin
        end
        8'hd7:
        begin
        end
        8'hd8:
        begin
        end
        8'hd9:
        begin
        end
        8'hda:
        begin
        end
        8'hdb:
        begin
        end
        8'hdc:
        begin
        end
        8'hdd:
        begin
        end
        8'hde:
        begin
        end
        8'hdf:
        begin
        end
        8'he0:
        begin
        end
        8'he1:
        begin
        end
        8'he2:
        begin
        end
        8'he3:
        begin
        end
        8'he4:
        begin
        end
        8'he5:
        begin
        end
        8'he6:
        begin
        end
        8'he7:
        begin
        end
        8'he8:
        begin
        end
        8'he9:
        begin
        end
        8'hea:
        begin
        end
        8'heb:
        begin
        end
        8'hec:
        begin
        end
        8'hed:
        begin
        end
        8'hee:
        begin
        end
        8'hef:
        begin
        end
        8'hf0:
        begin
        end
        8'hf1:
        begin
        end
        8'hf2:
        begin
        end
        8'hf3:
        begin
        end
        8'hf4:
        begin
        end
        8'hf5:
        begin
        end
        8'hf6:
        begin
        end
        8'hf7:
        begin
        end
        8'hf8:
        begin
        end
        8'hf9:
        begin
        end
        8'hfa:
        begin
        end
        8'hfb:
        begin
        end
        8'hfc:
        begin
        end
        8'hfd:
        begin
        end
        8'hfe:
        begin
        end
        8'hff:
        begin
        end
        endcase
    end
    assign \AES.rf.S4_4.out  = { \AES.rf.S4_4.k0 , \AES.rf.S4_4.k1 , \AES.rf.S4_4.k2 , \AES.rf.S4_4.k3  };
    assign \AES.rf.z0  = ( { \AES.rf.p00 , \AES.rf.p11 , \AES.rf.p22 , \AES.rf.p33  } ^ \AES.rf.k0  );
    assign \AES.rf.z1  = ( { \AES.rf.p10 , \AES.rf.p21 , \AES.rf.p32 , \AES.rf.p03  } ^ \AES.rf.k1  );
    assign \AES.rf.z2  = ( { \AES.rf.p20 , \AES.rf.p31 , \AES.rf.p02 , \AES.rf.p13  } ^ \AES.rf.k2  );
    assign \AES.rf.z3  = ( { \AES.rf.p30 , \AES.rf.p01 , \AES.rf.p12 , \AES.rf.p23  } ^ \AES.rf.k3  );
    always @ (  posedge \AES.rf.clk )
    begin
    end
endmodule 


