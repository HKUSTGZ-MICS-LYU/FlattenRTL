module wrapper #(
    parameter RTL__csr_regfile__f_reset_rsps__RTL__csr_regfile__guarded=32'd1,
    parameter RTL__stage1_f_reset_reqs__RTL__guarded=32'd1,
    parameter RTL__stage1_f_reset_rsps__RTL__guarded=32'd1,
    parameter RTL__stage2_f_reset_reqs__RTL__guarded=32'd1,
    parameter RTL__stage2_f_reset_rsps__RTL__guarded=32'd1,
    parameter RTL__stage3_f_reset_reqs__RTL__guarded=32'd1,
    parameter RTL__stage3_f_reset_rsps__RTL__guarded=32'd1,
parameter RTL__f_reset_reqs__RTL__width=32'd1,
parameter RTL__f_reset_reqs__RTL__guarded=32'd1,
parameter RTL__f_reset_rsps__RTL__width=32'd1,
parameter RTL__f_reset_rsps__RTL__guarded=32'd1,
parameter RTL__gpr_regfile__f_reset_rsps__RTL__gpr_regfile__guarded=32'd1,
parameter RTL__gpr_regfile__regfile__RTL__gpr_regfile__addr_width=32'd5,
parameter RTL__gpr_regfile__regfile__RTL__gpr_regfile__data_width=32'd32,
parameter RTL__gpr_regfile__regfile__RTL__gpr_regfile__lo=5'h0,
parameter RTL__gpr_regfile__regfile__RTL__gpr_regfile__hi=5'd31,
parameter RTL__near_mem__dcache__RTL__near_mem__dmem_not_imem=1'd1,
parameter RTL__near_mem__icache__RTL__near_mem__dmem_not_imem=1'd0,
parameter RTL__near_mem__dcache__f_fabric_write_reqs__RTL__near_mem__dcache__width=32'd99,
parameter RTL__near_mem__dcache__f_fabric_write_reqs__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__f_reset_reqs__RTL__near_mem__dcache__width=32'd1,
parameter RTL__near_mem__dcache__f_reset_reqs__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__f_reset_rsps__RTL__near_mem__dcache__width=32'd1,
parameter RTL__near_mem__dcache__f_reset_rsps__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__near_mem__dcache__width=32'd97,
parameter RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__near_mem__dcache__width=32'd71,
parameter RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__near_mem__dcache__width=32'd97,
parameter RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__near_mem__dcache__width=32'd73,
parameter RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__near_mem__dcache__width=32'd6,
parameter RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__near_mem__dcache__guarded=32'd1,
parameter RTL__near_mem__icache__f_fabric_write_reqs__RTL__near_mem__icache__width=32'd99,
parameter RTL__near_mem__icache__f_fabric_write_reqs__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__f_reset_reqs__RTL__near_mem__icache__width=32'd1,
parameter RTL__near_mem__icache__f_reset_reqs__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__f_reset_rsps__RTL__near_mem__icache__width=32'd1,
parameter RTL__near_mem__icache__f_reset_rsps__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__near_mem__icache__width=32'd97,
parameter RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__master_xactor_f_rd_data__RTL__near_mem__icache__width=32'd71,
parameter RTL__near_mem__icache__master_xactor_f_rd_data__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__near_mem__icache__width=32'd97,
parameter RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__master_xactor_f_wr_data__RTL__near_mem__icache__width=32'd73,
parameter RTL__near_mem__icache__master_xactor_f_wr_data__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__near_mem__icache__width=32'd6,
parameter RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__near_mem__icache__guarded=32'd1,
parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__RTL__near_mem__dcache__PIPELINED=1'd0,
parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__RTL__near_mem__dcache__ADDR_WIDTH=32'd7,
parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__RTL__near_mem__dcache__DATA_WIDTH=32'd23,
parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__RTL__near_mem__dcache__MEMSIZE=8'd128,
parameter RTL__near_mem__dcache__ram_word64_set__RTL__near_mem__dcache__PIPELINED=1'd0,
parameter RTL__near_mem__dcache__ram_word64_set__RTL__near_mem__dcache__ADDR_WIDTH=32'd9,
parameter RTL__near_mem__dcache__ram_word64_set__RTL__near_mem__dcache__DATA_WIDTH=32'd64,
parameter RTL__near_mem__dcache__ram_word64_set__RTL__near_mem__dcache__MEMSIZE=10'd512,
parameter RTL__near_mem__icache__ram_state_and_ctag_cset__RTL__near_mem__icache__PIPELINED=1'd0,
parameter RTL__near_mem__icache__ram_state_and_ctag_cset__RTL__near_mem__icache__ADDR_WIDTH=32'd7,
parameter RTL__near_mem__icache__ram_state_and_ctag_cset__RTL__near_mem__icache__DATA_WIDTH=32'd23,
parameter RTL__near_mem__icache__ram_state_and_ctag_cset__RTL__near_mem__icache__MEMSIZE=8'd128,
parameter RTL__near_mem__icache__ram_word64_set__RTL__near_mem__icache__PIPELINED=1'd0,
parameter RTL__near_mem__icache__ram_word64_set__RTL__near_mem__icache__ADDR_WIDTH=32'd9,
parameter RTL__near_mem__icache__ram_word64_set__RTL__near_mem__icache__DATA_WIDTH=32'd64,
parameter RTL__near_mem__icache__ram_word64_set__RTL__near_mem__icache__MEMSIZE=10'd512,
parameter RTL__near_mem__f_reset_rsps__RTL__near_mem__guarded=32'd1)(
__ILA_I_inst,
__ISSUE__,
__VLG_I_EN_hart0_server_reset_request_put,
__VLG_I_EN_hart0_server_reset_response_get,
__VLG_I_EN_set_verbosity,
__VLG_I_dmem_master_arready,
__VLG_I_dmem_master_awready,
__VLG_I_dmem_master_bid,
__VLG_I_dmem_master_bresp,
__VLG_I_dmem_master_bvalid,
__VLG_I_dmem_master_rdata,
__VLG_I_dmem_master_rid,
__VLG_I_dmem_master_rlast,
__VLG_I_dmem_master_rresp,
__VLG_I_dmem_master_rvalid,
__VLG_I_dmem_master_wready,
__VLG_I_hart0_server_reset_request_put,
__VLG_I_imem_master_arready,
__VLG_I_imem_master_awready,
__VLG_I_imem_master_bid,
__VLG_I_imem_master_bresp,
__VLG_I_imem_master_bvalid,
__VLG_I_imem_master_rdata,
__VLG_I_imem_master_rid,
__VLG_I_imem_master_rlast,
__VLG_I_imem_master_rresp,
__VLG_I_imem_master_rvalid,
__VLG_I_imem_master_wready,
__VLG_I_set_verbosity_logdelay,
__VLG_I_set_verbosity_verbosity,
____auxvar10__recorder_init__,
____auxvar11__recorder_init__,
____auxvar12__recorder_init__,
____auxvar13__recorder_init__,
____auxvar14__recorder_init__,
____auxvar15__recorder_init__,
____auxvar16__recorder_init__,
____auxvar17__recorder_init__,
____auxvar18__recorder_init__,
____auxvar19__recorder_init__,
____auxvar1__recorder_init__,
____auxvar20__recorder_init__,
____auxvar21__recorder_init__,
____auxvar22__recorder_init__,
____auxvar23__recorder_init__,
____auxvar24__recorder_init__,
____auxvar25__recorder_init__,
____auxvar26__recorder_init__,
____auxvar27__recorder_init__,
____auxvar28__recorder_init__,
____auxvar29__recorder_init__,
____auxvar2__recorder_init__,
____auxvar30__recorder_init__,
____auxvar31__recorder_init__,
____auxvar32__recorder_init__,
____auxvar33__recorder_init__,
____auxvar34__recorder_init__,
____auxvar35__recorder_init__,
____auxvar36__recorder_init__,
____auxvar37__recorder_init__,
____auxvar38__recorder_init__,
____auxvar3__recorder_init__,
____auxvar4__recorder_init__,
____auxvar5__recorder_init__,
____auxvar6__recorder_init__,
____auxvar7__recorder_init__,
____auxvar8__recorder_init__,
____auxvar9__recorder_init__,
clk,
dummy_reset,
rst,
RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__csr_regfile__DOT__rg_nmi,
RTL__DOT__csr_regfile__DOT__rg_state,
RTL__DOT__f_reset_reqs__DOT__empty_reg,
RTL__DOT__f_reset_reqs__DOT__full_reg,
RTL__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_,
RTL__DOT__near_mem$EN_dmem_req,
RTL__DOT__near_mem$dmem_exc,
RTL__DOT__near_mem$dmem_req_addr,
RTL__DOT__near_mem$dmem_req_f3,
RTL__DOT__near_mem$dmem_req_op,
RTL__DOT__near_mem$dmem_req_store_value,
RTL__DOT__near_mem$dmem_word64,
RTL__DOT__near_mem$imem_instr,
RTL__DOT__near_mem$imem_pc,
RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr,
RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa,
RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg,
RTL__DOT__rg_cur_priv,
RTL__DOT__rg_retiring$EN,
RTL__DOT__rg_run_on_reset,
RTL__DOT__rg_state,
RTL__DOT__rg_trap_instr,
RTL__DOT__s1_to_s2$D_IN,
RTL__DOT__s1_to_s2$EN,
RTL__DOT__s2_to_s3$D_IN,
RTL__DOT__s2_to_s3$EN,
RTL__DOT__s3_deq$D_IN,
RTL__DOT__s3_deq$EN,
RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg,
RTL__DOT__stage1_f_reset_reqs__DOT__full_reg,
RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg,
RTL__DOT__stage1_f_reset_rsps__DOT__full_reg,
RTL__DOT__stage1_rg_full,
RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg,
RTL__DOT__stage2_f_reset_reqs__DOT__full_reg,
RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg,
RTL__DOT__stage2_f_reset_rsps__DOT__full_reg,
RTL__DOT__stage2_rg_full,
RTL__DOT__stage2_rg_stage2,
RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg,
RTL__DOT__stage3_f_reset_reqs__DOT__full_reg,
RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg,
RTL__DOT__stage3_f_reset_rsps__DOT__full_reg,
RTL__DOT__stage3_rg_full,
__EDCOND__,
__IEND__,
__ILA_SO_load_addr,
__ILA_SO_load_data,
__ILA_SO_load_en,
__ILA_SO_load_size,
__ILA_SO_pc,
__ILA_SO_store_addr,
__ILA_SO_store_data,
__ILA_SO_store_en,
__ILA_SO_store_size,
__ILA_SO_x0,
__ILA_SO_x1,
__ILA_SO_x10,
__ILA_SO_x11,
__ILA_SO_x12,
__ILA_SO_x13,
__ILA_SO_x14,
__ILA_SO_x15,
__ILA_SO_x16,
__ILA_SO_x17,
__ILA_SO_x18,
__ILA_SO_x19,
__ILA_SO_x2,
__ILA_SO_x20,
__ILA_SO_x21,
__ILA_SO_x22,
__ILA_SO_x23,
__ILA_SO_x24,
__ILA_SO_x25,
__ILA_SO_x26,
__ILA_SO_x27,
__ILA_SO_x28,
__ILA_SO_x29,
__ILA_SO_x3,
__ILA_SO_x30,
__ILA_SO_x31,
__ILA_SO_x4,
__ILA_SO_x5,
__ILA_SO_x6,
__ILA_SO_x7,
__ILA_SO_x8,
__ILA_SO_x9,
__VLG_II_m_external_interrupt_req_set_not_clear,
__VLG_II_nmi_req_set_not_clear,
__VLG_II_s_external_interrupt_req_set_not_clear,
__VLG_II_software_interrupt_req_set_not_clear,
__VLG_II_timer_interrupt_req_set_not_clear,
__VLG_O_RDY_hart0_server_reset_request_put,
__VLG_O_RDY_hart0_server_reset_response_get,
__VLG_O_RDY_set_verbosity,
__VLG_O_dmem_master_araddr,
__VLG_O_dmem_master_arburst,
__VLG_O_dmem_master_arcache,
__VLG_O_dmem_master_arid,
__VLG_O_dmem_master_arlen,
__VLG_O_dmem_master_arlock,
__VLG_O_dmem_master_arprot,
__VLG_O_dmem_master_arqos,
__VLG_O_dmem_master_arregion,
__VLG_O_dmem_master_arsize,
__VLG_O_dmem_master_arvalid,
__VLG_O_dmem_master_awaddr,
__VLG_O_dmem_master_awburst,
__VLG_O_dmem_master_awcache,
__VLG_O_dmem_master_awid,
__VLG_O_dmem_master_awlen,
__VLG_O_dmem_master_awlock,
__VLG_O_dmem_master_awprot,
__VLG_O_dmem_master_awqos,
__VLG_O_dmem_master_awregion,
__VLG_O_dmem_master_awsize,
__VLG_O_dmem_master_awvalid,
__VLG_O_dmem_master_bready,
__VLG_O_dmem_master_rready,
__VLG_O_dmem_master_wdata,
__VLG_O_dmem_master_wlast,
__VLG_O_dmem_master_wstrb,
__VLG_O_dmem_master_wvalid,
__VLG_O_hart0_server_reset_response_get,
__VLG_O_imem_master_araddr,
__VLG_O_imem_master_arburst,
__VLG_O_imem_master_arcache,
__VLG_O_imem_master_arid,
__VLG_O_imem_master_arlen,
__VLG_O_imem_master_arlock,
__VLG_O_imem_master_arprot,
__VLG_O_imem_master_arqos,
__VLG_O_imem_master_arregion,
__VLG_O_imem_master_arsize,
__VLG_O_imem_master_arvalid,
__VLG_O_imem_master_awaddr,
__VLG_O_imem_master_awburst,
__VLG_O_imem_master_awcache,
__VLG_O_imem_master_awid,
__VLG_O_imem_master_awlen,
__VLG_O_imem_master_awlock,
__VLG_O_imem_master_awprot,
__VLG_O_imem_master_awqos,
__VLG_O_imem_master_awregion,
__VLG_O_imem_master_awsize,
__VLG_O_imem_master_awvalid,
__VLG_O_imem_master_bready,
__VLG_O_imem_master_rready,
__VLG_O_imem_master_wdata,
__VLG_O_imem_master_wlast,
__VLG_O_imem_master_wstrb,
__VLG_O_imem_master_wvalid,
__all_assert_wire__,
__all_assume_wire__,
__auxvar0__delay_d_0,
__sanitycheck_wire__,
end_of_pipeline,
input_map_assume___p0__,
invariant_assume__p10__,
invariant_assume__p11__,
invariant_assume__p12__,
invariant_assume__p13__,
invariant_assume__p14__,
invariant_assume__p15__,
invariant_assume__p16__,
invariant_assume__p17__,
invariant_assume__p18__,
invariant_assume__p19__,
invariant_assume__p1__,
invariant_assume__p20__,
invariant_assume__p21__,
invariant_assume__p22__,
invariant_assume__p23__,
invariant_assume__p24__,
invariant_assume__p25__,
invariant_assume__p26__,
invariant_assume__p27__,
invariant_assume__p28__,
invariant_assume__p29__,
invariant_assume__p2__,
invariant_assume__p30__,
invariant_assume__p31__,
invariant_assume__p32__,
invariant_assume__p3__,
invariant_assume__p4__,
invariant_assume__p5__,
invariant_assume__p6__,
invariant_assume__p7__,
invariant_assume__p8__,
invariant_assume__p9__,
issue_decode__p33__,
issue_valid__p34__,
mem_req_addr,
mem_req_en,
mem_req_funct3,
mem_req_op,
mem_req_rd_data,
mem_req_wd_data,
monitor_s1,
monitor_s1_already_enter_cond,
monitor_s1_already_exit_cond,
monitor_s2_enter_cond,
monitor_s2_exit_cond,
monitor_s3_enter_cond,
monitor_s3_exit_cond,
monitor_s4_enter_cond,
monitor_s4_exit_cond,
noreset__p35__,
post_value_holder__p36__,
post_value_holder__p37__,
post_value_holder__p38__,
post_value_holder__p39__,
post_value_holder__p40__,
post_value_holder__p41__,
post_value_holder__p42__,
post_value_holder__p43__,
post_value_holder__p44__,
post_value_holder__p45__,
post_value_holder__p46__,
post_value_holder__p47__,
post_value_holder__p48__,
post_value_holder__p49__,
post_value_holder__p50__,
post_value_holder__p51__,
post_value_holder__p52__,
post_value_holder__p53__,
post_value_holder__p54__,
post_value_holder__p55__,
post_value_holder__p56__,
post_value_holder__p57__,
post_value_holder__p58__,
post_value_holder__p59__,
post_value_holder__p60__,
post_value_holder__p61__,
post_value_holder__p62__,
post_value_holder__p63__,
post_value_holder__p64__,
post_value_holder__p65__,
post_value_holder__p66__,
post_value_holder__p67__,
post_value_holder__p68__,
post_value_holder__p69__,
post_value_holder__p70__,
post_value_holder__p71__,
post_value_holder__p72__,
post_value_holder__p73__,
post_value_holder_overly_constrained__p153__,
post_value_holder_overly_constrained__p154__,
post_value_holder_overly_constrained__p155__,
post_value_holder_overly_constrained__p156__,
post_value_holder_overly_constrained__p157__,
post_value_holder_overly_constrained__p158__,
post_value_holder_overly_constrained__p159__,
post_value_holder_overly_constrained__p160__,
post_value_holder_overly_constrained__p161__,
post_value_holder_overly_constrained__p162__,
post_value_holder_overly_constrained__p163__,
post_value_holder_overly_constrained__p164__,
post_value_holder_overly_constrained__p165__,
post_value_holder_overly_constrained__p166__,
post_value_holder_overly_constrained__p167__,
post_value_holder_overly_constrained__p168__,
post_value_holder_overly_constrained__p169__,
post_value_holder_overly_constrained__p170__,
post_value_holder_overly_constrained__p171__,
post_value_holder_overly_constrained__p172__,
post_value_holder_overly_constrained__p173__,
post_value_holder_overly_constrained__p174__,
post_value_holder_overly_constrained__p175__,
post_value_holder_overly_constrained__p176__,
post_value_holder_overly_constrained__p177__,
post_value_holder_overly_constrained__p178__,
post_value_holder_overly_constrained__p179__,
post_value_holder_overly_constrained__p180__,
post_value_holder_overly_constrained__p181__,
post_value_holder_overly_constrained__p182__,
post_value_holder_overly_constrained__p183__,
post_value_holder_overly_constrained__p184__,
post_value_holder_overly_constrained__p185__,
post_value_holder_overly_constrained__p186__,
post_value_holder_overly_constrained__p187__,
post_value_holder_overly_constrained__p188__,
post_value_holder_overly_constrained__p189__,
post_value_holder_overly_constrained__p190__,
post_value_holder_triggered__p191__,
post_value_holder_triggered__p192__,
post_value_holder_triggered__p193__,
post_value_holder_triggered__p194__,
post_value_holder_triggered__p195__,
post_value_holder_triggered__p196__,
post_value_holder_triggered__p197__,
post_value_holder_triggered__p198__,
post_value_holder_triggered__p199__,
post_value_holder_triggered__p200__,
post_value_holder_triggered__p201__,
post_value_holder_triggered__p202__,
post_value_holder_triggered__p203__,
post_value_holder_triggered__p204__,
post_value_holder_triggered__p205__,
post_value_holder_triggered__p206__,
post_value_holder_triggered__p207__,
post_value_holder_triggered__p208__,
post_value_holder_triggered__p209__,
post_value_holder_triggered__p210__,
post_value_holder_triggered__p211__,
post_value_holder_triggered__p212__,
post_value_holder_triggered__p213__,
post_value_holder_triggered__p214__,
post_value_holder_triggered__p215__,
post_value_holder_triggered__p216__,
post_value_holder_triggered__p217__,
post_value_holder_triggered__p218__,
post_value_holder_triggered__p219__,
post_value_holder_triggered__p220__,
post_value_holder_triggered__p221__,
post_value_holder_triggered__p222__,
post_value_holder_triggered__p223__,
post_value_holder_triggered__p224__,
post_value_holder_triggered__p225__,
post_value_holder_triggered__p226__,
post_value_holder_triggered__p227__,
post_value_holder_triggered__p228__,
rfassumptions__p74__,
rfassumptions__p75__,
rfassumptions__p76__,
s2_enter,
s2_exit,
s3_enter,
s3_exit,
s4_enter,
variable_map_assert__p118__,
variable_map_assert__p119__,
variable_map_assert__p120__,
variable_map_assert__p121__,
variable_map_assert__p122__,
variable_map_assert__p123__,
variable_map_assert__p124__,
variable_map_assert__p125__,
variable_map_assert__p126__,
variable_map_assert__p127__,
variable_map_assert__p128__,
variable_map_assert__p129__,
variable_map_assert__p130__,
variable_map_assert__p131__,
variable_map_assert__p132__,
variable_map_assert__p133__,
variable_map_assert__p134__,
variable_map_assert__p135__,
variable_map_assert__p136__,
variable_map_assert__p137__,
variable_map_assert__p138__,
variable_map_assert__p139__,
variable_map_assert__p140__,
variable_map_assert__p141__,
variable_map_assert__p142__,
variable_map_assert__p143__,
variable_map_assert__p144__,
variable_map_assert__p145__,
variable_map_assert__p146__,
variable_map_assert__p147__,
variable_map_assert__p148__,
variable_map_assert__p149__,
variable_map_assert__p150__,
variable_map_assert__p151__,
variable_map_assert__p152__,
variable_map_assume___p100__,
variable_map_assume___p101__,
variable_map_assume___p102__,
variable_map_assume___p103__,
variable_map_assume___p104__,
variable_map_assume___p105__,
variable_map_assume___p106__,
variable_map_assume___p107__,
variable_map_assume___p108__,
variable_map_assume___p109__,
variable_map_assume___p110__,
variable_map_assume___p111__,
variable_map_assume___p112__,
variable_map_assume___p113__,
variable_map_assume___p114__,
variable_map_assume___p115__,
variable_map_assume___p116__,
variable_map_assume___p117__,
variable_map_assume___p77__,
variable_map_assume___p78__,
variable_map_assume___p79__,
variable_map_assume___p80__,
variable_map_assume___p81__,
variable_map_assume___p82__,
variable_map_assume___p83__,
variable_map_assume___p84__,
variable_map_assume___p85__,
variable_map_assume___p86__,
variable_map_assume___p87__,
variable_map_assume___p88__,
variable_map_assume___p89__,
variable_map_assume___p90__,
variable_map_assume___p91__,
variable_map_assume___p92__,
variable_map_assume___p93__,
variable_map_assume___p94__,
variable_map_assume___p95__,
variable_map_assume___p96__,
variable_map_assume___p97__,
variable_map_assume___p98__,
variable_map_assume___p99__,
__CYCLE_CNT__,
__START__,
__STARTED__,
__ENDED__,
__2ndENDED__,
__RESETED__,
__auxvar10__recorder,
__auxvar10__recorder_sn_vhold,
__auxvar10__recorder_sn_condmet,
__auxvar11__recorder,
__auxvar11__recorder_sn_vhold,
__auxvar11__recorder_sn_condmet,
__auxvar12__recorder,
__auxvar12__recorder_sn_vhold,
__auxvar12__recorder_sn_condmet,
__auxvar13__recorder,
__auxvar13__recorder_sn_vhold,
__auxvar13__recorder_sn_condmet,
__auxvar14__recorder,
__auxvar14__recorder_sn_vhold,
__auxvar14__recorder_sn_condmet,
__auxvar15__recorder,
__auxvar15__recorder_sn_vhold,
__auxvar15__recorder_sn_condmet,
__auxvar16__recorder,
__auxvar16__recorder_sn_vhold,
__auxvar16__recorder_sn_condmet,
__auxvar17__recorder,
__auxvar17__recorder_sn_vhold,
__auxvar17__recorder_sn_condmet,
__auxvar18__recorder,
__auxvar18__recorder_sn_vhold,
__auxvar18__recorder_sn_condmet,
__auxvar19__recorder,
__auxvar19__recorder_sn_vhold,
__auxvar19__recorder_sn_condmet,
__auxvar1__recorder,
__auxvar1__recorder_sn_vhold,
__auxvar1__recorder_sn_condmet,
__auxvar20__recorder,
__auxvar20__recorder_sn_vhold,
__auxvar20__recorder_sn_condmet,
__auxvar21__recorder,
__auxvar21__recorder_sn_vhold,
__auxvar21__recorder_sn_condmet,
__auxvar22__recorder,
__auxvar22__recorder_sn_vhold,
__auxvar22__recorder_sn_condmet,
__auxvar23__recorder,
__auxvar23__recorder_sn_vhold,
__auxvar23__recorder_sn_condmet,
__auxvar24__recorder,
__auxvar24__recorder_sn_vhold,
__auxvar24__recorder_sn_condmet,
__auxvar25__recorder,
__auxvar25__recorder_sn_vhold,
__auxvar25__recorder_sn_condmet,
__auxvar26__recorder,
__auxvar26__recorder_sn_vhold,
__auxvar26__recorder_sn_condmet,
__auxvar27__recorder,
__auxvar27__recorder_sn_vhold,
__auxvar27__recorder_sn_condmet,
__auxvar28__recorder,
__auxvar28__recorder_sn_vhold,
__auxvar28__recorder_sn_condmet,
__auxvar29__recorder,
__auxvar29__recorder_sn_vhold,
__auxvar29__recorder_sn_condmet,
__auxvar2__recorder,
__auxvar2__recorder_sn_vhold,
__auxvar2__recorder_sn_condmet,
__auxvar30__recorder,
__auxvar30__recorder_sn_vhold,
__auxvar30__recorder_sn_condmet,
__auxvar31__recorder,
__auxvar31__recorder_sn_vhold,
__auxvar31__recorder_sn_condmet,
__auxvar32__recorder,
__auxvar32__recorder_sn_vhold,
__auxvar32__recorder_sn_condmet,
__auxvar33__recorder,
__auxvar33__recorder_sn_vhold,
__auxvar33__recorder_sn_condmet,
__auxvar34__recorder,
__auxvar34__recorder_sn_vhold,
__auxvar34__recorder_sn_condmet,
__auxvar35__recorder,
__auxvar35__recorder_sn_vhold,
__auxvar35__recorder_sn_condmet,
__auxvar36__recorder,
__auxvar36__recorder_sn_vhold,
__auxvar36__recorder_sn_condmet,
__auxvar37__recorder,
__auxvar37__recorder_sn_vhold,
__auxvar37__recorder_sn_condmet,
__auxvar38__recorder,
__auxvar38__recorder_sn_vhold,
__auxvar38__recorder_sn_condmet,
__auxvar3__recorder,
__auxvar3__recorder_sn_vhold,
__auxvar3__recorder_sn_condmet,
__auxvar4__recorder,
__auxvar4__recorder_sn_vhold,
__auxvar4__recorder_sn_condmet,
__auxvar5__recorder,
__auxvar5__recorder_sn_vhold,
__auxvar5__recorder_sn_condmet,
__auxvar6__recorder,
__auxvar6__recorder_sn_vhold,
__auxvar6__recorder_sn_condmet,
__auxvar7__recorder,
__auxvar7__recorder_sn_vhold,
__auxvar7__recorder_sn_condmet,
__auxvar8__recorder,
__auxvar8__recorder_sn_vhold,
__auxvar8__recorder_sn_condmet,
__auxvar9__recorder,
__auxvar9__recorder_sn_vhold,
__auxvar9__recorder_sn_condmet,
__auxvar0__delay_d_1,
monitor_s1_already,
monitor_s2,
monitor_s3,
monitor_s4
);
input     [31:0] __ILA_I_inst;
input            __ISSUE__;
input            __VLG_I_EN_hart0_server_reset_request_put;
input            __VLG_I_EN_hart0_server_reset_response_get;
input            __VLG_I_EN_set_verbosity;
input            __VLG_I_dmem_master_arready;
input            __VLG_I_dmem_master_awready;
input      [3:0] __VLG_I_dmem_master_bid;
input      [1:0] __VLG_I_dmem_master_bresp;
input            __VLG_I_dmem_master_bvalid;
input     [63:0] __VLG_I_dmem_master_rdata;
input      [3:0] __VLG_I_dmem_master_rid;
input            __VLG_I_dmem_master_rlast;
input      [1:0] __VLG_I_dmem_master_rresp;
input            __VLG_I_dmem_master_rvalid;
input            __VLG_I_dmem_master_wready;
input            __VLG_I_hart0_server_reset_request_put;
input            __VLG_I_imem_master_arready;
input            __VLG_I_imem_master_awready;
input      [3:0] __VLG_I_imem_master_bid;
input      [1:0] __VLG_I_imem_master_bresp;
input            __VLG_I_imem_master_bvalid;
input     [63:0] __VLG_I_imem_master_rdata;
input      [3:0] __VLG_I_imem_master_rid;
input            __VLG_I_imem_master_rlast;
input      [1:0] __VLG_I_imem_master_rresp;
input            __VLG_I_imem_master_rvalid;
input            __VLG_I_imem_master_wready;
input     [63:0] __VLG_I_set_verbosity_logdelay;
input      [3:0] __VLG_I_set_verbosity_verbosity;
input     [31:0] ____auxvar10__recorder_init__;
input     [31:0] ____auxvar11__recorder_init__;
input     [31:0] ____auxvar12__recorder_init__;
input     [31:0] ____auxvar13__recorder_init__;
input     [31:0] ____auxvar14__recorder_init__;
input     [31:0] ____auxvar15__recorder_init__;
input     [31:0] ____auxvar16__recorder_init__;
input     [31:0] ____auxvar17__recorder_init__;
input     [31:0] ____auxvar18__recorder_init__;
input     [31:0] ____auxvar19__recorder_init__;
input     [31:0] ____auxvar1__recorder_init__;
input     [31:0] ____auxvar20__recorder_init__;
input     [31:0] ____auxvar21__recorder_init__;
input     [31:0] ____auxvar22__recorder_init__;
input     [31:0] ____auxvar23__recorder_init__;
input     [31:0] ____auxvar24__recorder_init__;
input     [31:0] ____auxvar25__recorder_init__;
input     [31:0] ____auxvar26__recorder_init__;
input     [31:0] ____auxvar27__recorder_init__;
input     [31:0] ____auxvar28__recorder_init__;
input     [31:0] ____auxvar29__recorder_init__;
input     [31:0] ____auxvar2__recorder_init__;
input     [31:0] ____auxvar30__recorder_init__;
input     [31:0] ____auxvar31__recorder_init__;
input     [31:0] ____auxvar32__recorder_init__;
input     [31:0] ____auxvar33__recorder_init__;
input            ____auxvar34__recorder_init__;
input      [2:0] ____auxvar35__recorder_init__;
input            ____auxvar36__recorder_init__;
input     [31:0] ____auxvar37__recorder_init__;
input     [31:0] ____auxvar38__recorder_init__;
input     [31:0] ____auxvar3__recorder_init__;
input     [31:0] ____auxvar4__recorder_init__;
input     [31:0] ____auxvar5__recorder_init__;
input     [31:0] ____auxvar6__recorder_init__;
input     [31:0] ____auxvar7__recorder_init__;
input     [31:0] ____auxvar8__recorder_init__;
input     [31:0] ____auxvar9__recorder_init__;
input            clk;
input            dummy_reset;
input            rst;
output            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__csr_regfile__DOT__rg_nmi;
output            RTL__DOT__csr_regfile__DOT__rg_state;
output            RTL__DOT__f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__f_reset_reqs__DOT__full_reg;
output            RTL__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
output            RTL__DOT__near_mem$EN_dmem_req;
output            RTL__DOT__near_mem$dmem_exc;
output     [31:0] RTL__DOT__near_mem$dmem_req_addr;
output      [2:0] RTL__DOT__near_mem$dmem_req_f3;
output            RTL__DOT__near_mem$dmem_req_op;
output     [63:0] RTL__DOT__near_mem$dmem_req_store_value;
output     [63:0] RTL__DOT__near_mem$dmem_word64;
output     [31:0] RTL__DOT__near_mem$imem_instr;
output     [31:0] RTL__DOT__near_mem$imem_pc;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
output     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
output     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
output            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
output      [1:0] RTL__DOT__rg_cur_priv;
output            RTL__DOT__rg_retiring$EN;
output            RTL__DOT__rg_run_on_reset;
output      [3:0] RTL__DOT__rg_state;
output     [31:0] RTL__DOT__rg_trap_instr;
output            RTL__DOT__s1_to_s2$D_IN;
output            RTL__DOT__s1_to_s2$EN;
output            RTL__DOT__s2_to_s3$D_IN;
output            RTL__DOT__s2_to_s3$EN;
output            RTL__DOT__s3_deq$D_IN;
output            RTL__DOT__s3_deq$EN;
output            RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
output            RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
output            RTL__DOT__stage1_rg_full;
output            RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
output            RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
output            RTL__DOT__stage2_rg_full;
output    [168:0] RTL__DOT__stage2_rg_stage2;
output            RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
output            RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
output            RTL__DOT__stage3_rg_full;
output            __EDCOND__;
output            __IEND__;
output     [31:0] __ILA_SO_load_addr;
output     [31:0] __ILA_SO_load_data;
output            __ILA_SO_load_en;
output      [2:0] __ILA_SO_load_size;
output     [31:0] __ILA_SO_pc;
output     [31:0] __ILA_SO_store_addr;
output     [31:0] __ILA_SO_store_data;
output            __ILA_SO_store_en;
output      [2:0] __ILA_SO_store_size;
output     [31:0] __ILA_SO_x0;
output     [31:0] __ILA_SO_x1;
output     [31:0] __ILA_SO_x10;
output     [31:0] __ILA_SO_x11;
output     [31:0] __ILA_SO_x12;
output     [31:0] __ILA_SO_x13;
output     [31:0] __ILA_SO_x14;
output     [31:0] __ILA_SO_x15;
output     [31:0] __ILA_SO_x16;
output     [31:0] __ILA_SO_x17;
output     [31:0] __ILA_SO_x18;
output     [31:0] __ILA_SO_x19;
output     [31:0] __ILA_SO_x2;
output     [31:0] __ILA_SO_x20;
output     [31:0] __ILA_SO_x21;
output     [31:0] __ILA_SO_x22;
output     [31:0] __ILA_SO_x23;
output     [31:0] __ILA_SO_x24;
output     [31:0] __ILA_SO_x25;
output     [31:0] __ILA_SO_x26;
output     [31:0] __ILA_SO_x27;
output     [31:0] __ILA_SO_x28;
output     [31:0] __ILA_SO_x29;
output     [31:0] __ILA_SO_x3;
output     [31:0] __ILA_SO_x30;
output     [31:0] __ILA_SO_x31;
output     [31:0] __ILA_SO_x4;
output     [31:0] __ILA_SO_x5;
output     [31:0] __ILA_SO_x6;
output     [31:0] __ILA_SO_x7;
output     [31:0] __ILA_SO_x8;
output     [31:0] __ILA_SO_x9;
output            __VLG_II_m_external_interrupt_req_set_not_clear;
output            __VLG_II_nmi_req_set_not_clear;
output            __VLG_II_s_external_interrupt_req_set_not_clear;
output            __VLG_II_software_interrupt_req_set_not_clear;
output            __VLG_II_timer_interrupt_req_set_not_clear;
output            __VLG_O_RDY_hart0_server_reset_request_put;
output            __VLG_O_RDY_hart0_server_reset_response_get;
output            __VLG_O_RDY_set_verbosity;
output     [63:0] __VLG_O_dmem_master_araddr;
output      [1:0] __VLG_O_dmem_master_arburst;
output      [3:0] __VLG_O_dmem_master_arcache;
output      [3:0] __VLG_O_dmem_master_arid;
output      [7:0] __VLG_O_dmem_master_arlen;
output            __VLG_O_dmem_master_arlock;
output      [2:0] __VLG_O_dmem_master_arprot;
output      [3:0] __VLG_O_dmem_master_arqos;
output      [3:0] __VLG_O_dmem_master_arregion;
output      [2:0] __VLG_O_dmem_master_arsize;
output            __VLG_O_dmem_master_arvalid;
output     [63:0] __VLG_O_dmem_master_awaddr;
output      [1:0] __VLG_O_dmem_master_awburst;
output      [3:0] __VLG_O_dmem_master_awcache;
output      [3:0] __VLG_O_dmem_master_awid;
output      [7:0] __VLG_O_dmem_master_awlen;
output            __VLG_O_dmem_master_awlock;
output      [2:0] __VLG_O_dmem_master_awprot;
output      [3:0] __VLG_O_dmem_master_awqos;
output      [3:0] __VLG_O_dmem_master_awregion;
output      [2:0] __VLG_O_dmem_master_awsize;
output            __VLG_O_dmem_master_awvalid;
output            __VLG_O_dmem_master_bready;
output            __VLG_O_dmem_master_rready;
output     [63:0] __VLG_O_dmem_master_wdata;
output            __VLG_O_dmem_master_wlast;
output      [7:0] __VLG_O_dmem_master_wstrb;
output            __VLG_O_dmem_master_wvalid;
output            __VLG_O_hart0_server_reset_response_get;
output     [63:0] __VLG_O_imem_master_araddr;
output      [1:0] __VLG_O_imem_master_arburst;
output      [3:0] __VLG_O_imem_master_arcache;
output      [3:0] __VLG_O_imem_master_arid;
output      [7:0] __VLG_O_imem_master_arlen;
output            __VLG_O_imem_master_arlock;
output      [2:0] __VLG_O_imem_master_arprot;
output      [3:0] __VLG_O_imem_master_arqos;
output      [3:0] __VLG_O_imem_master_arregion;
output      [2:0] __VLG_O_imem_master_arsize;
output            __VLG_O_imem_master_arvalid;
output     [63:0] __VLG_O_imem_master_awaddr;
output      [1:0] __VLG_O_imem_master_awburst;
output      [3:0] __VLG_O_imem_master_awcache;
output      [3:0] __VLG_O_imem_master_awid;
output      [7:0] __VLG_O_imem_master_awlen;
output            __VLG_O_imem_master_awlock;
output      [2:0] __VLG_O_imem_master_awprot;
output      [3:0] __VLG_O_imem_master_awqos;
output      [3:0] __VLG_O_imem_master_awregion;
output      [2:0] __VLG_O_imem_master_awsize;
output            __VLG_O_imem_master_awvalid;
output            __VLG_O_imem_master_bready;
output            __VLG_O_imem_master_rready;
output     [63:0] __VLG_O_imem_master_wdata;
output            __VLG_O_imem_master_wlast;
output      [7:0] __VLG_O_imem_master_wstrb;
output            __VLG_O_imem_master_wvalid;
output            __all_assert_wire__;
output            __all_assume_wire__;
output            __auxvar0__delay_d_0;
output            __sanitycheck_wire__;
output            end_of_pipeline;
output            input_map_assume___p0__;
output            invariant_assume__p10__;
output            invariant_assume__p11__;
output            invariant_assume__p12__;
output            invariant_assume__p13__;
output            invariant_assume__p14__;
output            invariant_assume__p15__;
output            invariant_assume__p16__;
output            invariant_assume__p17__;
output            invariant_assume__p18__;
output            invariant_assume__p19__;
output            invariant_assume__p1__;
output            invariant_assume__p20__;
output            invariant_assume__p21__;
output            invariant_assume__p22__;
output            invariant_assume__p23__;
output            invariant_assume__p24__;
output            invariant_assume__p25__;
output            invariant_assume__p26__;
output            invariant_assume__p27__;
output            invariant_assume__p28__;
output            invariant_assume__p29__;
output            invariant_assume__p2__;
output            invariant_assume__p30__;
output            invariant_assume__p31__;
output            invariant_assume__p32__;
output            invariant_assume__p3__;
output            invariant_assume__p4__;
output            invariant_assume__p5__;
output            invariant_assume__p6__;
output            invariant_assume__p7__;
output            invariant_assume__p8__;
output            invariant_assume__p9__;
output            issue_decode__p33__;
output            issue_valid__p34__;
output     [31:0] mem_req_addr;
output            mem_req_en;
output      [2:0] mem_req_funct3;
output            mem_req_op;
output     [31:0] mem_req_rd_data;
output     [31:0] mem_req_wd_data;
output            monitor_s1;
output            monitor_s1_already_enter_cond;
output            monitor_s1_already_exit_cond;
output            monitor_s2_enter_cond;
output            monitor_s2_exit_cond;
output            monitor_s3_enter_cond;
output            monitor_s3_exit_cond;
output            monitor_s4_enter_cond;
output            monitor_s4_exit_cond;
output            noreset__p35__;
output            post_value_holder__p36__;
output            post_value_holder__p37__;
output            post_value_holder__p38__;
output            post_value_holder__p39__;
output            post_value_holder__p40__;
output            post_value_holder__p41__;
output            post_value_holder__p42__;
output            post_value_holder__p43__;
output            post_value_holder__p44__;
output            post_value_holder__p45__;
output            post_value_holder__p46__;
output            post_value_holder__p47__;
output            post_value_holder__p48__;
output            post_value_holder__p49__;
output            post_value_holder__p50__;
output            post_value_holder__p51__;
output            post_value_holder__p52__;
output            post_value_holder__p53__;
output            post_value_holder__p54__;
output            post_value_holder__p55__;
output            post_value_holder__p56__;
output            post_value_holder__p57__;
output            post_value_holder__p58__;
output            post_value_holder__p59__;
output            post_value_holder__p60__;
output            post_value_holder__p61__;
output            post_value_holder__p62__;
output            post_value_holder__p63__;
output            post_value_holder__p64__;
output            post_value_holder__p65__;
output            post_value_holder__p66__;
output            post_value_holder__p67__;
output            post_value_holder__p68__;
output            post_value_holder__p69__;
output            post_value_holder__p70__;
output            post_value_holder__p71__;
output            post_value_holder__p72__;
output            post_value_holder__p73__;
output            post_value_holder_overly_constrained__p153__;
output            post_value_holder_overly_constrained__p154__;
output            post_value_holder_overly_constrained__p155__;
output            post_value_holder_overly_constrained__p156__;
output            post_value_holder_overly_constrained__p157__;
output            post_value_holder_overly_constrained__p158__;
output            post_value_holder_overly_constrained__p159__;
output            post_value_holder_overly_constrained__p160__;
output            post_value_holder_overly_constrained__p161__;
output            post_value_holder_overly_constrained__p162__;
output            post_value_holder_overly_constrained__p163__;
output            post_value_holder_overly_constrained__p164__;
output            post_value_holder_overly_constrained__p165__;
output            post_value_holder_overly_constrained__p166__;
output            post_value_holder_overly_constrained__p167__;
output            post_value_holder_overly_constrained__p168__;
output            post_value_holder_overly_constrained__p169__;
output            post_value_holder_overly_constrained__p170__;
output            post_value_holder_overly_constrained__p171__;
output            post_value_holder_overly_constrained__p172__;
output            post_value_holder_overly_constrained__p173__;
output            post_value_holder_overly_constrained__p174__;
output            post_value_holder_overly_constrained__p175__;
output            post_value_holder_overly_constrained__p176__;
output            post_value_holder_overly_constrained__p177__;
output            post_value_holder_overly_constrained__p178__;
output            post_value_holder_overly_constrained__p179__;
output            post_value_holder_overly_constrained__p180__;
output            post_value_holder_overly_constrained__p181__;
output            post_value_holder_overly_constrained__p182__;
output            post_value_holder_overly_constrained__p183__;
output            post_value_holder_overly_constrained__p184__;
output            post_value_holder_overly_constrained__p185__;
output            post_value_holder_overly_constrained__p186__;
output            post_value_holder_overly_constrained__p187__;
output            post_value_holder_overly_constrained__p188__;
output            post_value_holder_overly_constrained__p189__;
output            post_value_holder_overly_constrained__p190__;
output            post_value_holder_triggered__p191__;
output            post_value_holder_triggered__p192__;
output            post_value_holder_triggered__p193__;
output            post_value_holder_triggered__p194__;
output            post_value_holder_triggered__p195__;
output            post_value_holder_triggered__p196__;
output            post_value_holder_triggered__p197__;
output            post_value_holder_triggered__p198__;
output            post_value_holder_triggered__p199__;
output            post_value_holder_triggered__p200__;
output            post_value_holder_triggered__p201__;
output            post_value_holder_triggered__p202__;
output            post_value_holder_triggered__p203__;
output            post_value_holder_triggered__p204__;
output            post_value_holder_triggered__p205__;
output            post_value_holder_triggered__p206__;
output            post_value_holder_triggered__p207__;
output            post_value_holder_triggered__p208__;
output            post_value_holder_triggered__p209__;
output            post_value_holder_triggered__p210__;
output            post_value_holder_triggered__p211__;
output            post_value_holder_triggered__p212__;
output            post_value_holder_triggered__p213__;
output            post_value_holder_triggered__p214__;
output            post_value_holder_triggered__p215__;
output            post_value_holder_triggered__p216__;
output            post_value_holder_triggered__p217__;
output            post_value_holder_triggered__p218__;
output            post_value_holder_triggered__p219__;
output            post_value_holder_triggered__p220__;
output            post_value_holder_triggered__p221__;
output            post_value_holder_triggered__p222__;
output            post_value_holder_triggered__p223__;
output            post_value_holder_triggered__p224__;
output            post_value_holder_triggered__p225__;
output            post_value_holder_triggered__p226__;
output            post_value_holder_triggered__p227__;
output            post_value_holder_triggered__p228__;
output            rfassumptions__p74__;
output            rfassumptions__p75__;
output            rfassumptions__p76__;
output            s2_enter;
output            s2_exit;
output            s3_enter;
output            s3_exit;
output            s4_enter;
output            variable_map_assert__p118__;
output            variable_map_assert__p119__;
output            variable_map_assert__p120__;
output            variable_map_assert__p121__;
output            variable_map_assert__p122__;
output            variable_map_assert__p123__;
output            variable_map_assert__p124__;
output            variable_map_assert__p125__;
output            variable_map_assert__p126__;
output            variable_map_assert__p127__;
output            variable_map_assert__p128__;
output            variable_map_assert__p129__;
output            variable_map_assert__p130__;
output            variable_map_assert__p131__;
output            variable_map_assert__p132__;
output            variable_map_assert__p133__;
output            variable_map_assert__p134__;
output            variable_map_assert__p135__;
output            variable_map_assert__p136__;
output            variable_map_assert__p137__;
output            variable_map_assert__p138__;
output            variable_map_assert__p139__;
output            variable_map_assert__p140__;
output            variable_map_assert__p141__;
output            variable_map_assert__p142__;
output            variable_map_assert__p143__;
output            variable_map_assert__p144__;
output            variable_map_assert__p145__;
output            variable_map_assert__p146__;
output            variable_map_assert__p147__;
output            variable_map_assert__p148__;
output            variable_map_assert__p149__;
output            variable_map_assert__p150__;
output            variable_map_assert__p151__;
output            variable_map_assert__p152__;
output            variable_map_assume___p100__;
output            variable_map_assume___p101__;
output            variable_map_assume___p102__;
output            variable_map_assume___p103__;
output            variable_map_assume___p104__;
output            variable_map_assume___p105__;
output            variable_map_assume___p106__;
output            variable_map_assume___p107__;
output            variable_map_assume___p108__;
output            variable_map_assume___p109__;
output            variable_map_assume___p110__;
output            variable_map_assume___p111__;
output            variable_map_assume___p112__;
output            variable_map_assume___p113__;
output            variable_map_assume___p114__;
output            variable_map_assume___p115__;
output            variable_map_assume___p116__;
output            variable_map_assume___p117__;
output            variable_map_assume___p77__;
output            variable_map_assume___p78__;
output            variable_map_assume___p79__;
output            variable_map_assume___p80__;
output            variable_map_assume___p81__;
output            variable_map_assume___p82__;
output            variable_map_assume___p83__;
output            variable_map_assume___p84__;
output            variable_map_assume___p85__;
output            variable_map_assume___p86__;
output            variable_map_assume___p87__;
output            variable_map_assume___p88__;
output            variable_map_assume___p89__;
output            variable_map_assume___p90__;
output            variable_map_assume___p91__;
output            variable_map_assume___p92__;
output            variable_map_assume___p93__;
output            variable_map_assume___p94__;
output            variable_map_assume___p95__;
output            variable_map_assume___p96__;
output            variable_map_assume___p97__;
output            variable_map_assume___p98__;
output            variable_map_assume___p99__;
output reg      [7:0] __CYCLE_CNT__;
output reg            __START__;
output reg            __STARTED__;
output reg            __ENDED__;
output reg            __2ndENDED__;
output reg            __RESETED__;
output reg     [31:0] __auxvar10__recorder;
output reg     [31:0] __auxvar10__recorder_sn_vhold;
output reg            __auxvar10__recorder_sn_condmet;
output reg     [31:0] __auxvar11__recorder;
output reg     [31:0] __auxvar11__recorder_sn_vhold;
output reg            __auxvar11__recorder_sn_condmet;
output reg     [31:0] __auxvar12__recorder;
output reg     [31:0] __auxvar12__recorder_sn_vhold;
output reg            __auxvar12__recorder_sn_condmet;
output reg     [31:0] __auxvar13__recorder;
output reg     [31:0] __auxvar13__recorder_sn_vhold;
output reg            __auxvar13__recorder_sn_condmet;
output reg     [31:0] __auxvar14__recorder;
output reg     [31:0] __auxvar14__recorder_sn_vhold;
output reg            __auxvar14__recorder_sn_condmet;
output reg     [31:0] __auxvar15__recorder;
output reg     [31:0] __auxvar15__recorder_sn_vhold;
output reg            __auxvar15__recorder_sn_condmet;
output reg     [31:0] __auxvar16__recorder;
output reg     [31:0] __auxvar16__recorder_sn_vhold;
output reg            __auxvar16__recorder_sn_condmet;
output reg     [31:0] __auxvar17__recorder;
output reg     [31:0] __auxvar17__recorder_sn_vhold;
output reg            __auxvar17__recorder_sn_condmet;
output reg     [31:0] __auxvar18__recorder;
output reg     [31:0] __auxvar18__recorder_sn_vhold;
output reg            __auxvar18__recorder_sn_condmet;
output reg     [31:0] __auxvar19__recorder;
output reg     [31:0] __auxvar19__recorder_sn_vhold;
output reg            __auxvar19__recorder_sn_condmet;
output reg     [31:0] __auxvar1__recorder;
output reg     [31:0] __auxvar1__recorder_sn_vhold;
output reg            __auxvar1__recorder_sn_condmet;
output reg     [31:0] __auxvar20__recorder;
output reg     [31:0] __auxvar20__recorder_sn_vhold;
output reg            __auxvar20__recorder_sn_condmet;
output reg     [31:0] __auxvar21__recorder;
output reg     [31:0] __auxvar21__recorder_sn_vhold;
output reg            __auxvar21__recorder_sn_condmet;
output reg     [31:0] __auxvar22__recorder;
output reg     [31:0] __auxvar22__recorder_sn_vhold;
output reg            __auxvar22__recorder_sn_condmet;
output reg     [31:0] __auxvar23__recorder;
output reg     [31:0] __auxvar23__recorder_sn_vhold;
output reg            __auxvar23__recorder_sn_condmet;
output reg     [31:0] __auxvar24__recorder;
output reg     [31:0] __auxvar24__recorder_sn_vhold;
output reg            __auxvar24__recorder_sn_condmet;
output reg     [31:0] __auxvar25__recorder;
output reg     [31:0] __auxvar25__recorder_sn_vhold;
output reg            __auxvar25__recorder_sn_condmet;
output reg     [31:0] __auxvar26__recorder;
output reg     [31:0] __auxvar26__recorder_sn_vhold;
output reg            __auxvar26__recorder_sn_condmet;
output reg     [31:0] __auxvar27__recorder;
output reg     [31:0] __auxvar27__recorder_sn_vhold;
output reg            __auxvar27__recorder_sn_condmet;
output reg     [31:0] __auxvar28__recorder;
output reg     [31:0] __auxvar28__recorder_sn_vhold;
output reg            __auxvar28__recorder_sn_condmet;
output reg     [31:0] __auxvar29__recorder;
output reg     [31:0] __auxvar29__recorder_sn_vhold;
output reg            __auxvar29__recorder_sn_condmet;
output reg     [31:0] __auxvar2__recorder;
output reg     [31:0] __auxvar2__recorder_sn_vhold;
output reg            __auxvar2__recorder_sn_condmet;
output reg     [31:0] __auxvar30__recorder;
output reg     [31:0] __auxvar30__recorder_sn_vhold;
output reg            __auxvar30__recorder_sn_condmet;
output reg     [31:0] __auxvar31__recorder;
output reg     [31:0] __auxvar31__recorder_sn_vhold;
output reg            __auxvar31__recorder_sn_condmet;
output reg     [31:0] __auxvar32__recorder;
output reg     [31:0] __auxvar32__recorder_sn_vhold;
output reg            __auxvar32__recorder_sn_condmet;
output reg     [31:0] __auxvar33__recorder;
output reg     [31:0] __auxvar33__recorder_sn_vhold;
output reg            __auxvar33__recorder_sn_condmet;
output reg            __auxvar34__recorder;
output reg            __auxvar34__recorder_sn_vhold;
output reg            __auxvar34__recorder_sn_condmet;
output reg      [2:0] __auxvar35__recorder;
output reg      [2:0] __auxvar35__recorder_sn_vhold;
output reg            __auxvar35__recorder_sn_condmet;
output reg            __auxvar36__recorder;
output reg            __auxvar36__recorder_sn_vhold;
output reg            __auxvar36__recorder_sn_condmet;
output reg     [31:0] __auxvar37__recorder;
output reg     [31:0] __auxvar37__recorder_sn_vhold;
output reg            __auxvar37__recorder_sn_condmet;
output reg     [31:0] __auxvar38__recorder;
output reg     [31:0] __auxvar38__recorder_sn_vhold;
output reg            __auxvar38__recorder_sn_condmet;
output reg     [31:0] __auxvar3__recorder;
output reg     [31:0] __auxvar3__recorder_sn_vhold;
output reg            __auxvar3__recorder_sn_condmet;
output reg     [31:0] __auxvar4__recorder;
output reg     [31:0] __auxvar4__recorder_sn_vhold;
output reg            __auxvar4__recorder_sn_condmet;
output reg     [31:0] __auxvar5__recorder;
output reg     [31:0] __auxvar5__recorder_sn_vhold;
output reg            __auxvar5__recorder_sn_condmet;
output reg     [31:0] __auxvar6__recorder;
output reg     [31:0] __auxvar6__recorder_sn_vhold;
output reg            __auxvar6__recorder_sn_condmet;
output reg     [31:0] __auxvar7__recorder;
output reg     [31:0] __auxvar7__recorder_sn_vhold;
output reg            __auxvar7__recorder_sn_condmet;
output reg     [31:0] __auxvar8__recorder;
output reg     [31:0] __auxvar8__recorder_sn_vhold;
output reg            __auxvar8__recorder_sn_condmet;
output reg     [31:0] __auxvar9__recorder;
output reg     [31:0] __auxvar9__recorder_sn_vhold;
output reg            __auxvar9__recorder_sn_condmet;
output reg            __auxvar0__delay_d_1;
output reg            monitor_s1_already;
output reg            monitor_s2;
output reg            monitor_s3;
output reg            monitor_s4;
(* keep *) wire            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__csr_regfile__DOT__rg_nmi;
(* keep *) wire            RTL__DOT__csr_regfile__DOT__rg_state;
(* keep *) wire            RTL__DOT__f_reset_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__f_reset_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
(* keep *) wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
(* keep *) wire            RTL__DOT__near_mem$EN_dmem_req;
(* keep *) wire            RTL__DOT__near_mem$dmem_exc;
(* keep *) wire     [31:0] RTL__DOT__near_mem$dmem_req_addr;
(* keep *) wire      [2:0] RTL__DOT__near_mem$dmem_req_f3;
(* keep *) wire            RTL__DOT__near_mem$dmem_req_op;
(* keep *) wire     [63:0] RTL__DOT__near_mem$dmem_req_store_value;
(* keep *) wire     [63:0] RTL__DOT__near_mem$dmem_word64;
(* keep *) wire     [31:0] RTL__DOT__near_mem$imem_instr;
(* keep *) wire     [31:0] RTL__DOT__near_mem$imem_pc;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
(* keep *) wire     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
(* keep *) wire     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
(* keep *) wire            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
(* keep *) wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
(* keep *) wire      [1:0] RTL__DOT__rg_cur_priv;
(* keep *) wire            RTL__DOT__rg_retiring$EN;
(* keep *) wire            RTL__DOT__rg_run_on_reset;
(* keep *) wire      [3:0] RTL__DOT__rg_state;
(* keep *) wire     [31:0] RTL__DOT__rg_trap_instr;
(* keep *) wire            RTL__DOT__s1_to_s2$D_IN;
(* keep *) wire            RTL__DOT__s1_to_s2$EN;
(* keep *) wire            RTL__DOT__s2_to_s3$D_IN;
(* keep *) wire            RTL__DOT__s2_to_s3$EN;
(* keep *) wire            RTL__DOT__s3_deq$D_IN;
(* keep *) wire            RTL__DOT__s3_deq$EN;
(* keep *) wire            RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__stage1_rg_full;
(* keep *) wire            RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__stage2_rg_full;
(* keep *) wire    [168:0] RTL__DOT__stage2_rg_stage2;
(* keep *) wire            RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
(* keep *) wire            RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
(* keep *) wire            RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
(* keep *) wire            RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
(* keep *) wire            RTL__DOT__stage3_rg_full;
wire            __2ndIEND__;
(* keep *) wire            __EDCOND__;
(* keep *) wire            __IEND__;
(* keep *) wire     [31:0] __ILA_I_inst;
(* keep *) wire     [31:0] __ILA_SO_load_addr;
(* keep *) wire     [31:0] __ILA_SO_load_data;
(* keep *) wire            __ILA_SO_load_en;
(* keep *) wire      [2:0] __ILA_SO_load_size;
(* keep *) wire     [31:0] __ILA_SO_pc;
(* keep *) wire     [31:0] __ILA_SO_store_addr;
(* keep *) wire     [31:0] __ILA_SO_store_data;
(* keep *) wire            __ILA_SO_store_en;
(* keep *) wire      [2:0] __ILA_SO_store_size;
(* keep *) wire     [31:0] __ILA_SO_x0;
(* keep *) wire     [31:0] __ILA_SO_x1;
(* keep *) wire     [31:0] __ILA_SO_x10;
(* keep *) wire     [31:0] __ILA_SO_x11;
(* keep *) wire     [31:0] __ILA_SO_x12;
(* keep *) wire     [31:0] __ILA_SO_x13;
(* keep *) wire     [31:0] __ILA_SO_x14;
(* keep *) wire     [31:0] __ILA_SO_x15;
(* keep *) wire     [31:0] __ILA_SO_x16;
(* keep *) wire     [31:0] __ILA_SO_x17;
(* keep *) wire     [31:0] __ILA_SO_x18;
(* keep *) wire     [31:0] __ILA_SO_x19;
(* keep *) wire     [31:0] __ILA_SO_x2;
(* keep *) wire     [31:0] __ILA_SO_x20;
(* keep *) wire     [31:0] __ILA_SO_x21;
(* keep *) wire     [31:0] __ILA_SO_x22;
(* keep *) wire     [31:0] __ILA_SO_x23;
(* keep *) wire     [31:0] __ILA_SO_x24;
(* keep *) wire     [31:0] __ILA_SO_x25;
(* keep *) wire     [31:0] __ILA_SO_x26;
(* keep *) wire     [31:0] __ILA_SO_x27;
(* keep *) wire     [31:0] __ILA_SO_x28;
(* keep *) wire     [31:0] __ILA_SO_x29;
(* keep *) wire     [31:0] __ILA_SO_x3;
(* keep *) wire     [31:0] __ILA_SO_x30;
(* keep *) wire     [31:0] __ILA_SO_x31;
(* keep *) wire     [31:0] __ILA_SO_x4;
(* keep *) wire     [31:0] __ILA_SO_x5;
(* keep *) wire     [31:0] __ILA_SO_x6;
(* keep *) wire     [31:0] __ILA_SO_x7;
(* keep *) wire     [31:0] __ILA_SO_x8;
(* keep *) wire     [31:0] __ILA_SO_x9;
(* keep *) wire            __ILA_riscv_decode_of_ADD__;
(* keep *) wire            __ILA_riscv_valid__;
(* keep *) wire            __ISSUE__;
(* keep *) wire            __VLG_II_m_external_interrupt_req_set_not_clear;
(* keep *) wire            __VLG_II_nmi_req_set_not_clear;
(* keep *) wire            __VLG_II_s_external_interrupt_req_set_not_clear;
(* keep *) wire            __VLG_II_software_interrupt_req_set_not_clear;
(* keep *) wire            __VLG_II_timer_interrupt_req_set_not_clear;
(* keep *) wire            __VLG_I_EN_hart0_server_reset_request_put;
(* keep *) wire            __VLG_I_EN_hart0_server_reset_response_get;
(* keep *) wire            __VLG_I_EN_set_verbosity;
(* keep *) wire            __VLG_I_dmem_master_arready;
(* keep *) wire            __VLG_I_dmem_master_awready;
(* keep *) wire      [3:0] __VLG_I_dmem_master_bid;
(* keep *) wire      [1:0] __VLG_I_dmem_master_bresp;
(* keep *) wire            __VLG_I_dmem_master_bvalid;
(* keep *) wire     [63:0] __VLG_I_dmem_master_rdata;
(* keep *) wire      [3:0] __VLG_I_dmem_master_rid;
(* keep *) wire            __VLG_I_dmem_master_rlast;
(* keep *) wire      [1:0] __VLG_I_dmem_master_rresp;
(* keep *) wire            __VLG_I_dmem_master_rvalid;
(* keep *) wire            __VLG_I_dmem_master_wready;
(* keep *) wire            __VLG_I_hart0_server_reset_request_put;
(* keep *) wire            __VLG_I_imem_master_arready;
(* keep *) wire            __VLG_I_imem_master_awready;
(* keep *) wire      [3:0] __VLG_I_imem_master_bid;
(* keep *) wire      [1:0] __VLG_I_imem_master_bresp;
(* keep *) wire            __VLG_I_imem_master_bvalid;
(* keep *) wire     [63:0] __VLG_I_imem_master_rdata;
(* keep *) wire      [3:0] __VLG_I_imem_master_rid;
(* keep *) wire            __VLG_I_imem_master_rlast;
(* keep *) wire      [1:0] __VLG_I_imem_master_rresp;
(* keep *) wire            __VLG_I_imem_master_rvalid;
(* keep *) wire            __VLG_I_imem_master_wready;
(* keep *) wire     [63:0] __VLG_I_set_verbosity_logdelay;
(* keep *) wire      [3:0] __VLG_I_set_verbosity_verbosity;
(* keep *) wire            __VLG_O_RDY_hart0_server_reset_request_put;
(* keep *) wire            __VLG_O_RDY_hart0_server_reset_response_get;
(* keep *) wire            __VLG_O_RDY_set_verbosity;
(* keep *) wire     [63:0] __VLG_O_dmem_master_araddr;
(* keep *) wire      [1:0] __VLG_O_dmem_master_arburst;
(* keep *) wire      [3:0] __VLG_O_dmem_master_arcache;
(* keep *) wire      [3:0] __VLG_O_dmem_master_arid;
(* keep *) wire      [7:0] __VLG_O_dmem_master_arlen;
(* keep *) wire            __VLG_O_dmem_master_arlock;
(* keep *) wire      [2:0] __VLG_O_dmem_master_arprot;
(* keep *) wire      [3:0] __VLG_O_dmem_master_arqos;
(* keep *) wire      [3:0] __VLG_O_dmem_master_arregion;
(* keep *) wire      [2:0] __VLG_O_dmem_master_arsize;
(* keep *) wire            __VLG_O_dmem_master_arvalid;
(* keep *) wire     [63:0] __VLG_O_dmem_master_awaddr;
(* keep *) wire      [1:0] __VLG_O_dmem_master_awburst;
(* keep *) wire      [3:0] __VLG_O_dmem_master_awcache;
(* keep *) wire      [3:0] __VLG_O_dmem_master_awid;
(* keep *) wire      [7:0] __VLG_O_dmem_master_awlen;
(* keep *) wire            __VLG_O_dmem_master_awlock;
(* keep *) wire      [2:0] __VLG_O_dmem_master_awprot;
(* keep *) wire      [3:0] __VLG_O_dmem_master_awqos;
(* keep *) wire      [3:0] __VLG_O_dmem_master_awregion;
(* keep *) wire      [2:0] __VLG_O_dmem_master_awsize;
(* keep *) wire            __VLG_O_dmem_master_awvalid;
(* keep *) wire            __VLG_O_dmem_master_bready;
(* keep *) wire            __VLG_O_dmem_master_rready;
(* keep *) wire     [63:0] __VLG_O_dmem_master_wdata;
(* keep *) wire            __VLG_O_dmem_master_wlast;
(* keep *) wire      [7:0] __VLG_O_dmem_master_wstrb;
(* keep *) wire            __VLG_O_dmem_master_wvalid;
(* keep *) wire            __VLG_O_hart0_server_reset_response_get;
(* keep *) wire     [63:0] __VLG_O_imem_master_araddr;
(* keep *) wire      [1:0] __VLG_O_imem_master_arburst;
(* keep *) wire      [3:0] __VLG_O_imem_master_arcache;
(* keep *) wire      [3:0] __VLG_O_imem_master_arid;
(* keep *) wire      [7:0] __VLG_O_imem_master_arlen;
(* keep *) wire            __VLG_O_imem_master_arlock;
(* keep *) wire      [2:0] __VLG_O_imem_master_arprot;
(* keep *) wire      [3:0] __VLG_O_imem_master_arqos;
(* keep *) wire      [3:0] __VLG_O_imem_master_arregion;
(* keep *) wire      [2:0] __VLG_O_imem_master_arsize;
(* keep *) wire            __VLG_O_imem_master_arvalid;
(* keep *) wire     [63:0] __VLG_O_imem_master_awaddr;
(* keep *) wire      [1:0] __VLG_O_imem_master_awburst;
(* keep *) wire      [3:0] __VLG_O_imem_master_awcache;
(* keep *) wire      [3:0] __VLG_O_imem_master_awid;
(* keep *) wire      [7:0] __VLG_O_imem_master_awlen;
(* keep *) wire            __VLG_O_imem_master_awlock;
(* keep *) wire      [2:0] __VLG_O_imem_master_awprot;
(* keep *) wire      [3:0] __VLG_O_imem_master_awqos;
(* keep *) wire      [3:0] __VLG_O_imem_master_awregion;
(* keep *) wire      [2:0] __VLG_O_imem_master_awsize;
(* keep *) wire            __VLG_O_imem_master_awvalid;
(* keep *) wire            __VLG_O_imem_master_bready;
(* keep *) wire            __VLG_O_imem_master_rready;
(* keep *) wire     [63:0] __VLG_O_imem_master_wdata;
(* keep *) wire            __VLG_O_imem_master_wlast;
(* keep *) wire      [7:0] __VLG_O_imem_master_wstrb;
(* keep *) wire            __VLG_O_imem_master_wvalid;
wire     [31:0] ____auxvar10__recorder_init__;
wire     [31:0] ____auxvar11__recorder_init__;
wire     [31:0] ____auxvar12__recorder_init__;
wire     [31:0] ____auxvar13__recorder_init__;
wire     [31:0] ____auxvar14__recorder_init__;
wire     [31:0] ____auxvar15__recorder_init__;
wire     [31:0] ____auxvar16__recorder_init__;
wire     [31:0] ____auxvar17__recorder_init__;
wire     [31:0] ____auxvar18__recorder_init__;
wire     [31:0] ____auxvar19__recorder_init__;
wire     [31:0] ____auxvar1__recorder_init__;
wire     [31:0] ____auxvar20__recorder_init__;
wire     [31:0] ____auxvar21__recorder_init__;
wire     [31:0] ____auxvar22__recorder_init__;
wire     [31:0] ____auxvar23__recorder_init__;
wire     [31:0] ____auxvar24__recorder_init__;
wire     [31:0] ____auxvar25__recorder_init__;
wire     [31:0] ____auxvar26__recorder_init__;
wire     [31:0] ____auxvar27__recorder_init__;
wire     [31:0] ____auxvar28__recorder_init__;
wire     [31:0] ____auxvar29__recorder_init__;
wire     [31:0] ____auxvar2__recorder_init__;
wire     [31:0] ____auxvar30__recorder_init__;
wire     [31:0] ____auxvar31__recorder_init__;
wire     [31:0] ____auxvar32__recorder_init__;
wire     [31:0] ____auxvar33__recorder_init__;
wire            ____auxvar34__recorder_init__;
wire      [2:0] ____auxvar35__recorder_init__;
wire            ____auxvar36__recorder_init__;
wire     [31:0] ____auxvar37__recorder_init__;
wire     [31:0] ____auxvar38__recorder_init__;
wire     [31:0] ____auxvar3__recorder_init__;
wire     [31:0] ____auxvar4__recorder_init__;
wire     [31:0] ____auxvar5__recorder_init__;
wire     [31:0] ____auxvar6__recorder_init__;
wire     [31:0] ____auxvar7__recorder_init__;
wire     [31:0] ____auxvar8__recorder_init__;
wire     [31:0] ____auxvar9__recorder_init__;
(* keep *) wire            __all_assert_wire__;
(* keep *) wire            __all_assume_wire__;
wire            __auxvar0__delay;
(* keep *) wire            __auxvar0__delay_d_0;
wire            __auxvar10__recorder_sn_cond;
wire     [31:0] __auxvar10__recorder_sn_value;
wire            __auxvar11__recorder_sn_cond;
wire     [31:0] __auxvar11__recorder_sn_value;
wire            __auxvar12__recorder_sn_cond;
wire     [31:0] __auxvar12__recorder_sn_value;
wire            __auxvar13__recorder_sn_cond;
wire     [31:0] __auxvar13__recorder_sn_value;
wire            __auxvar14__recorder_sn_cond;
wire     [31:0] __auxvar14__recorder_sn_value;
wire            __auxvar15__recorder_sn_cond;
wire     [31:0] __auxvar15__recorder_sn_value;
wire            __auxvar16__recorder_sn_cond;
wire     [31:0] __auxvar16__recorder_sn_value;
wire            __auxvar17__recorder_sn_cond;
wire     [31:0] __auxvar17__recorder_sn_value;
wire            __auxvar18__recorder_sn_cond;
wire     [31:0] __auxvar18__recorder_sn_value;
wire            __auxvar19__recorder_sn_cond;
wire     [31:0] __auxvar19__recorder_sn_value;
wire            __auxvar1__recorder_sn_cond;
wire     [31:0] __auxvar1__recorder_sn_value;
wire            __auxvar20__recorder_sn_cond;
wire     [31:0] __auxvar20__recorder_sn_value;
wire            __auxvar21__recorder_sn_cond;
wire     [31:0] __auxvar21__recorder_sn_value;
wire            __auxvar22__recorder_sn_cond;
wire     [31:0] __auxvar22__recorder_sn_value;
wire            __auxvar23__recorder_sn_cond;
wire     [31:0] __auxvar23__recorder_sn_value;
wire            __auxvar24__recorder_sn_cond;
wire     [31:0] __auxvar24__recorder_sn_value;
wire            __auxvar25__recorder_sn_cond;
wire     [31:0] __auxvar25__recorder_sn_value;
wire            __auxvar26__recorder_sn_cond;
wire     [31:0] __auxvar26__recorder_sn_value;
wire            __auxvar27__recorder_sn_cond;
wire     [31:0] __auxvar27__recorder_sn_value;
wire            __auxvar28__recorder_sn_cond;
wire     [31:0] __auxvar28__recorder_sn_value;
wire            __auxvar29__recorder_sn_cond;
wire     [31:0] __auxvar29__recorder_sn_value;
wire            __auxvar2__recorder_sn_cond;
wire     [31:0] __auxvar2__recorder_sn_value;
wire            __auxvar30__recorder_sn_cond;
wire     [31:0] __auxvar30__recorder_sn_value;
wire            __auxvar31__recorder_sn_cond;
wire     [31:0] __auxvar31__recorder_sn_value;
wire            __auxvar32__recorder_sn_cond;
wire     [31:0] __auxvar32__recorder_sn_value;
wire            __auxvar33__recorder_sn_cond;
wire     [31:0] __auxvar33__recorder_sn_value;
wire            __auxvar34__recorder_sn_cond;
wire            __auxvar34__recorder_sn_value;
wire            __auxvar35__recorder_sn_cond;
wire      [2:0] __auxvar35__recorder_sn_value;
wire            __auxvar36__recorder_sn_cond;
wire            __auxvar36__recorder_sn_value;
wire            __auxvar37__recorder_sn_cond;
wire     [31:0] __auxvar37__recorder_sn_value;
wire            __auxvar38__recorder_sn_cond;
wire     [31:0] __auxvar38__recorder_sn_value;
wire            __auxvar3__recorder_sn_cond;
wire     [31:0] __auxvar3__recorder_sn_value;
wire            __auxvar4__recorder_sn_cond;
wire     [31:0] __auxvar4__recorder_sn_value;
wire            __auxvar5__recorder_sn_cond;
wire     [31:0] __auxvar5__recorder_sn_value;
wire            __auxvar6__recorder_sn_cond;
wire     [31:0] __auxvar6__recorder_sn_value;
wire            __auxvar7__recorder_sn_cond;
wire     [31:0] __auxvar7__recorder_sn_value;
wire            __auxvar8__recorder_sn_cond;
wire     [31:0] __auxvar8__recorder_sn_value;
wire            __auxvar9__recorder_sn_cond;
wire     [31:0] __auxvar9__recorder_sn_value;
(* keep *) wire            __sanitycheck_wire__;
wire            clk;
(* keep *) wire            dummy_reset;
wire            end_of_pipeline;
wire            input_map_assume___p0__;
wire            invariant_assume__p10__;
wire            invariant_assume__p11__;
wire            invariant_assume__p12__;
wire            invariant_assume__p13__;
wire            invariant_assume__p14__;
wire            invariant_assume__p15__;
wire            invariant_assume__p16__;
wire            invariant_assume__p17__;
wire            invariant_assume__p18__;
wire            invariant_assume__p19__;
wire            invariant_assume__p1__;
wire            invariant_assume__p20__;
wire            invariant_assume__p21__;
wire            invariant_assume__p22__;
wire            invariant_assume__p23__;
wire            invariant_assume__p24__;
wire            invariant_assume__p25__;
wire            invariant_assume__p26__;
wire            invariant_assume__p27__;
wire            invariant_assume__p28__;
wire            invariant_assume__p29__;
wire            invariant_assume__p2__;
wire            invariant_assume__p30__;
wire            invariant_assume__p31__;
wire            invariant_assume__p32__;
wire            invariant_assume__p3__;
wire            invariant_assume__p4__;
wire            invariant_assume__p5__;
wire            invariant_assume__p6__;
wire            invariant_assume__p7__;
wire            invariant_assume__p8__;
wire            invariant_assume__p9__;
wire            issue_decode__p33__;
wire            issue_valid__p34__;
(* keep *) wire     [31:0] mem_req_addr;
(* keep *) wire            mem_req_en;
(* keep *) wire      [2:0] mem_req_funct3;
(* keep *) wire            mem_req_op;
(* keep *) wire     [31:0] mem_req_rd_data;
(* keep *) wire     [31:0] mem_req_wd_data;
wire            monitor_s1;
(* keep *) wire            monitor_s1_already_enter_cond;
(* keep *) wire            monitor_s1_already_exit_cond;
(* keep *) wire            monitor_s2_enter_cond;
(* keep *) wire            monitor_s2_exit_cond;
(* keep *) wire            monitor_s3_enter_cond;
(* keep *) wire            monitor_s3_exit_cond;
(* keep *) wire            monitor_s4_enter_cond;
(* keep *) wire            monitor_s4_exit_cond;
wire            noreset__p35__;
wire            post_value_holder__p36__;
wire            post_value_holder__p37__;
wire            post_value_holder__p38__;
wire            post_value_holder__p39__;
wire            post_value_holder__p40__;
wire            post_value_holder__p41__;
wire            post_value_holder__p42__;
wire            post_value_holder__p43__;
wire            post_value_holder__p44__;
wire            post_value_holder__p45__;
wire            post_value_holder__p46__;
wire            post_value_holder__p47__;
wire            post_value_holder__p48__;
wire            post_value_holder__p49__;
wire            post_value_holder__p50__;
wire            post_value_holder__p51__;
wire            post_value_holder__p52__;
wire            post_value_holder__p53__;
wire            post_value_holder__p54__;
wire            post_value_holder__p55__;
wire            post_value_holder__p56__;
wire            post_value_holder__p57__;
wire            post_value_holder__p58__;
wire            post_value_holder__p59__;
wire            post_value_holder__p60__;
wire            post_value_holder__p61__;
wire            post_value_holder__p62__;
wire            post_value_holder__p63__;
wire            post_value_holder__p64__;
wire            post_value_holder__p65__;
wire            post_value_holder__p66__;
wire            post_value_holder__p67__;
wire            post_value_holder__p68__;
wire            post_value_holder__p69__;
wire            post_value_holder__p70__;
wire            post_value_holder__p71__;
wire            post_value_holder__p72__;
wire            post_value_holder__p73__;
wire            post_value_holder_overly_constrained__p153__;
wire            post_value_holder_overly_constrained__p154__;
wire            post_value_holder_overly_constrained__p155__;
wire            post_value_holder_overly_constrained__p156__;
wire            post_value_holder_overly_constrained__p157__;
wire            post_value_holder_overly_constrained__p158__;
wire            post_value_holder_overly_constrained__p159__;
wire            post_value_holder_overly_constrained__p160__;
wire            post_value_holder_overly_constrained__p161__;
wire            post_value_holder_overly_constrained__p162__;
wire            post_value_holder_overly_constrained__p163__;
wire            post_value_holder_overly_constrained__p164__;
wire            post_value_holder_overly_constrained__p165__;
wire            post_value_holder_overly_constrained__p166__;
wire            post_value_holder_overly_constrained__p167__;
wire            post_value_holder_overly_constrained__p168__;
wire            post_value_holder_overly_constrained__p169__;
wire            post_value_holder_overly_constrained__p170__;
wire            post_value_holder_overly_constrained__p171__;
wire            post_value_holder_overly_constrained__p172__;
wire            post_value_holder_overly_constrained__p173__;
wire            post_value_holder_overly_constrained__p174__;
wire            post_value_holder_overly_constrained__p175__;
wire            post_value_holder_overly_constrained__p176__;
wire            post_value_holder_overly_constrained__p177__;
wire            post_value_holder_overly_constrained__p178__;
wire            post_value_holder_overly_constrained__p179__;
wire            post_value_holder_overly_constrained__p180__;
wire            post_value_holder_overly_constrained__p181__;
wire            post_value_holder_overly_constrained__p182__;
wire            post_value_holder_overly_constrained__p183__;
wire            post_value_holder_overly_constrained__p184__;
wire            post_value_holder_overly_constrained__p185__;
wire            post_value_holder_overly_constrained__p186__;
wire            post_value_holder_overly_constrained__p187__;
wire            post_value_holder_overly_constrained__p188__;
wire            post_value_holder_overly_constrained__p189__;
wire            post_value_holder_overly_constrained__p190__;
wire            post_value_holder_triggered__p191__;
wire            post_value_holder_triggered__p192__;
wire            post_value_holder_triggered__p193__;
wire            post_value_holder_triggered__p194__;
wire            post_value_holder_triggered__p195__;
wire            post_value_holder_triggered__p196__;
wire            post_value_holder_triggered__p197__;
wire            post_value_holder_triggered__p198__;
wire            post_value_holder_triggered__p199__;
wire            post_value_holder_triggered__p200__;
wire            post_value_holder_triggered__p201__;
wire            post_value_holder_triggered__p202__;
wire            post_value_holder_triggered__p203__;
wire            post_value_holder_triggered__p204__;
wire            post_value_holder_triggered__p205__;
wire            post_value_holder_triggered__p206__;
wire            post_value_holder_triggered__p207__;
wire            post_value_holder_triggered__p208__;
wire            post_value_holder_triggered__p209__;
wire            post_value_holder_triggered__p210__;
wire            post_value_holder_triggered__p211__;
wire            post_value_holder_triggered__p212__;
wire            post_value_holder_triggered__p213__;
wire            post_value_holder_triggered__p214__;
wire            post_value_holder_triggered__p215__;
wire            post_value_holder_triggered__p216__;
wire            post_value_holder_triggered__p217__;
wire            post_value_holder_triggered__p218__;
wire            post_value_holder_triggered__p219__;
wire            post_value_holder_triggered__p220__;
wire            post_value_holder_triggered__p221__;
wire            post_value_holder_triggered__p222__;
wire            post_value_holder_triggered__p223__;
wire            post_value_holder_triggered__p224__;
wire            post_value_holder_triggered__p225__;
wire            post_value_holder_triggered__p226__;
wire            post_value_holder_triggered__p227__;
wire            post_value_holder_triggered__p228__;
wire            rfassumptions__p74__;
wire            rfassumptions__p75__;
wire            rfassumptions__p76__;
wire            rst;
wire            s2_enter;
wire            s2_exit;
wire            s3_enter;
wire            s3_exit;
wire            s4_enter;
wire            variable_map_assert__p118__;
wire            variable_map_assert__p119__;
wire            variable_map_assert__p120__;
wire            variable_map_assert__p121__;
wire            variable_map_assert__p122__;
wire            variable_map_assert__p123__;
wire            variable_map_assert__p124__;
wire            variable_map_assert__p125__;
wire            variable_map_assert__p126__;
wire            variable_map_assert__p127__;
wire            variable_map_assert__p128__;
wire            variable_map_assert__p129__;
wire            variable_map_assert__p130__;
wire            variable_map_assert__p131__;
wire            variable_map_assert__p132__;
wire            variable_map_assert__p133__;
wire            variable_map_assert__p134__;
wire            variable_map_assert__p135__;
wire            variable_map_assert__p136__;
wire            variable_map_assert__p137__;
wire            variable_map_assert__p138__;
wire            variable_map_assert__p139__;
wire            variable_map_assert__p140__;
wire            variable_map_assert__p141__;
wire            variable_map_assert__p142__;
wire            variable_map_assert__p143__;
wire            variable_map_assert__p144__;
wire            variable_map_assert__p145__;
wire            variable_map_assert__p146__;
wire            variable_map_assert__p147__;
wire            variable_map_assert__p148__;
wire            variable_map_assert__p149__;
wire            variable_map_assert__p150__;
wire            variable_map_assert__p151__;
wire            variable_map_assert__p152__;
wire            variable_map_assume___p100__;
wire            variable_map_assume___p101__;
wire            variable_map_assume___p102__;
wire            variable_map_assume___p103__;
wire            variable_map_assume___p104__;
wire            variable_map_assume___p105__;
wire            variable_map_assume___p106__;
wire            variable_map_assume___p107__;
wire            variable_map_assume___p108__;
wire            variable_map_assume___p109__;
wire            variable_map_assume___p110__;
wire            variable_map_assume___p111__;
wire            variable_map_assume___p112__;
wire            variable_map_assume___p113__;
wire            variable_map_assume___p114__;
wire            variable_map_assume___p115__;
wire            variable_map_assume___p116__;
wire            variable_map_assume___p117__;
wire            variable_map_assume___p77__;
wire            variable_map_assume___p78__;
wire            variable_map_assume___p79__;
wire            variable_map_assume___p80__;
wire            variable_map_assume___p81__;
wire            variable_map_assume___p82__;
wire            variable_map_assume___p83__;
wire            variable_map_assume___p84__;
wire            variable_map_assume___p85__;
wire            variable_map_assume___p86__;
wire            variable_map_assume___p87__;
wire            variable_map_assume___p88__;
wire            variable_map_assume___p89__;
wire            variable_map_assume___p90__;
wire            variable_map_assume___p91__;
wire            variable_map_assume___p92__;
wire            variable_map_assume___p93__;
wire            variable_map_assume___p94__;
wire            variable_map_assume___p95__;
wire            variable_map_assume___p96__;
wire            variable_map_assume___p97__;
wire            variable_map_assume___p98__;
wire            variable_map_assume___p99__;
always @(posedge clk) begin
if (rst) __CYCLE_CNT__ <= 0;
else if ( ( __START__ || __STARTED__ ) &&  __CYCLE_CNT__ < 137) __CYCLE_CNT__ <= __CYCLE_CNT__ + 1;
end
always @(posedge clk) begin
if (__ISSUE__ && !__START__ && !__STARTED__) __START__ <= 1;
else if (__START__ || __STARTED__) __START__ <= 0;
end
always @(posedge clk) begin
if (rst) __STARTED__ <= 0;
else if (__START__) __STARTED__ <= 1;
end
always @(posedge clk) begin
if (rst) __ENDED__ <= 0;
else if (__IEND__) __ENDED__ <= 1;
end
always @(posedge clk) begin
if (rst) __2ndENDED__ <= 1'b0;
else if (__ENDED__ && __EDCOND__ && ~__2ndENDED__)  __2ndENDED__ <= 1'b1; end
assign __2ndIEND__ = __ENDED__ && __EDCOND__ && ~__2ndENDED__ ;
always @(posedge clk) begin
if (rst) __RESETED__ <= 1;
end
assign __auxvar0__delay = __auxvar0__delay_d_1 ;
assign monitor_s1_already_exit_cond = 1'b0 ;
assign monitor_s4_exit_cond = 1'b0 ;
    wire ILA____START__;
    wire ILA__clk;
    wire[31:0] ILA__inst;
    wire ILA__rst;
    wire ILA____ILA_riscv_decode_of_ADD__;
    wire ILA____ILA_riscv_valid__;
    reg[31:0] ILA__pc;
    reg ILA__load_en;
    reg[31:0] ILA__load_addr;
    reg[2:0] ILA__load_size;
    reg[31:0] ILA__load_data;
    reg ILA__store_en;
    reg[31:0] ILA__store_addr;
    reg[2:0] ILA__store_size;
    reg[31:0] ILA__store_data;
    reg[31:0] ILA__x0;
    reg[31:0] ILA__x1;
    reg[31:0] ILA__x2;
    reg[31:0] ILA__x3;
    reg[31:0] ILA__x4;
    reg[31:0] ILA__x5;
    reg[31:0] ILA__x6;
    reg[31:0] ILA__x7;
    reg[31:0] ILA__x8;
    reg[31:0] ILA__x9;
    reg[31:0] ILA__x10;
    reg[31:0] ILA__x11;
    reg[31:0] ILA__x12;
    reg[31:0] ILA__x13;
    reg[31:0] ILA__x14;
    reg[31:0] ILA__x15;
    reg[31:0] ILA__x16;
    reg[31:0] ILA__x17;
    reg[31:0] ILA__x18;
    reg[31:0] ILA__x19;
    reg[31:0] ILA__x20;
    reg[31:0] ILA__x21;
    reg[31:0] ILA__x22;
    reg[31:0] ILA__x23;
    reg[31:0] ILA__x24;
    reg[31:0] ILA__x25;
    reg[31:0] ILA__x26;
    reg[31:0] ILA__x27;
    reg[31:0] ILA__x28;
    reg[31:0] ILA__x29;
    reg[31:0] ILA__x30;
    reg[31:0] ILA__x31;
    reg[7:0] ILA____COUNTER_start__n11;

    wire ILA____ILA_riscv_decode_of_ADD__ ; 
    wire ILA____ILA_riscv_valid__ ; 
    wire ILA____START__ ; 
    wire ILA__bv_1_0_n14 ; 
    wire[31:0] ILA__bv_32_0_n15 ; 
    wire[31:0] ILA__bv_32_4_n12 ; 
    wire[2:0] ILA__bv_3_0_n4 ; 
    wire[4:0] ILA__bv_5_10_n62 ; 
    wire[4:0] ILA__bv_5_11_n60 ; 
    wire[4:0] ILA__bv_5_12_n58 ; 
    wire[4:0] ILA__bv_5_13_n56 ; 
    wire[4:0] ILA__bv_5_14_n54 ; 
    wire[4:0] ILA__bv_5_15_n52 ; 
    wire[4:0] ILA__bv_5_16_n50 ; 
    wire[4:0] ILA__bv_5_17_n48 ; 
    wire[4:0] ILA__bv_5_18_n46 ; 
    wire[4:0] ILA__bv_5_19_n44 ; 
    wire[4:0] ILA__bv_5_1_n17 ; 
    wire[4:0] ILA__bv_5_20_n42 ; 
    wire[4:0] ILA__bv_5_21_n40 ; 
    wire[4:0] ILA__bv_5_22_n38 ; 
    wire[4:0] ILA__bv_5_23_n36 ; 
    wire[4:0] ILA__bv_5_24_n34 ; 
    wire[4:0] ILA__bv_5_25_n32 ; 
    wire[4:0] ILA__bv_5_26_n30 ; 
    wire[4:0] ILA__bv_5_27_n28 ; 
    wire[4:0] ILA__bv_5_28_n26 ; 
    wire[4:0] ILA__bv_5_29_n24 ; 
    wire[4:0] ILA__bv_5_2_n78 ; 
    wire[4:0] ILA__bv_5_30_n22 ; 
    wire[4:0] ILA__bv_5_31_n20 ; 
    wire[4:0] ILA__bv_5_3_n76 ; 
    wire[4:0] ILA__bv_5_4_n74 ; 
    wire[4:0] ILA__bv_5_5_n72 ; 
    wire[4:0] ILA__bv_5_6_n70 ; 
    wire[4:0] ILA__bv_5_7_n68 ; 
    wire[4:0] ILA__bv_5_8_n66 ; 
    wire[4:0] ILA__bv_5_9_n64 ; 
    wire[6:0] ILA__bv_7_0_n8 ; 
    wire[6:0] ILA__bv_7_51_n1 ; 
    wire ILA__clk ; 
    wire[31:0] ILA__inst ; (* ILA__keep *)
    wire[31:0] ILA__load_addr_randinit ; (* ILA__keep *)
    wire[31:0] ILA__load_data_randinit ; (* ILA__keep *)
    wire ILA__load_en_randinit ; (* ILA__keep *)
    wire[2:0] ILA__load_size_randinit ; 
    wire[6:0] ILA__n0 ; 
    wire ILA__n10 ; 
    wire[31:0] ILA__n100 ; 
    wire[31:0] ILA__n101 ; 
    wire[31:0] ILA__n102 ; 
    wire[31:0] ILA__n103 ; 
    wire[31:0] ILA__n104 ; 
    wire[31:0] ILA__n105 ; 
    wire[31:0] ILA__n106 ; 
    wire[31:0] ILA__n107 ; 
    wire[31:0] ILA__n108 ; 
    wire[31:0] ILA__n109 ; 
    wire[31:0] ILA__n110 ; 
    wire[31:0] ILA__n111 ; 
    wire[4:0] ILA__n112 ; 
    wire ILA__n113 ; 
    wire ILA__n114 ; 
    wire ILA__n115 ; 
    wire ILA__n116 ; 
    wire ILA__n117 ; 
    wire ILA__n118 ; 
    wire ILA__n119 ; 
    wire ILA__n120 ; 
    wire ILA__n121 ; 
    wire ILA__n122 ; 
    wire ILA__n123 ; 
    wire ILA__n124 ; 
    wire ILA__n125 ; 
    wire ILA__n126 ; 
    wire ILA__n127 ; 
    wire ILA__n128 ; 
    wire ILA__n129 ; 
    wire[31:0] ILA__n13 ; 
    wire ILA__n130 ; 
    wire ILA__n131 ; 
    wire ILA__n132 ; 
    wire ILA__n133 ; 
    wire ILA__n134 ; 
    wire ILA__n135 ; 
    wire ILA__n136 ; 
    wire ILA__n137 ; 
    wire ILA__n138 ; 
    wire ILA__n139 ; 
    wire ILA__n140 ; 
    wire ILA__n141 ; 
    wire ILA__n142 ; 
    wire ILA__n143 ; 
    wire[31:0] ILA__n144 ; 
    wire[31:0] ILA__n145 ; 
    wire[31:0] ILA__n146 ; 
    wire[31:0] ILA__n147 ; 
    wire[31:0] ILA__n148 ; 
    wire[31:0] ILA__n149 ; 
    wire[31:0] ILA__n150 ; 
    wire[31:0] ILA__n151 ; 
    wire[31:0] ILA__n152 ; 
    wire[31:0] ILA__n153 ; 
    wire[31:0] ILA__n154 ; 
    wire[31:0] ILA__n155 ; 
    wire[31:0] ILA__n156 ; 
    wire[31:0] ILA__n157 ; 
    wire[31:0] ILA__n158 ; 
    wire[31:0] ILA__n159 ; 
    wire[4:0] ILA__n16 ; 
    wire[31:0] ILA__n160 ; 
    wire[31:0] ILA__n161 ; 
    wire[31:0] ILA__n162 ; 
    wire[31:0] ILA__n163 ; 
    wire[31:0] ILA__n164 ; 
    wire[31:0] ILA__n165 ; 
    wire[31:0] ILA__n166 ; 
    wire[31:0] ILA__n167 ; 
    wire[31:0] ILA__n168 ; 
    wire[31:0] ILA__n169 ; 
    wire[31:0] ILA__n170 ; 
    wire[31:0] ILA__n171 ; 
    wire[31:0] ILA__n172 ; 
    wire[31:0] ILA__n173 ; 
    wire[31:0] ILA__n174 ; 
    wire[31:0] ILA__n175 ; 
    wire[31:0] ILA__n176 ; 
    wire ILA__n177 ; 
    wire[31:0] ILA__n178 ; 
    wire ILA__n179 ; 
    wire ILA__n18 ; 
    wire[31:0] ILA__n180 ; 
    wire ILA__n181 ; 
    wire[31:0] ILA__n182 ; 
    wire ILA__n183 ; 
    wire[31:0] ILA__n184 ; 
    wire ILA__n185 ; 
    wire[31:0] ILA__n186 ; 
    wire ILA__n187 ; 
    wire[31:0] ILA__n188 ; 
    wire ILA__n189 ; 
    wire[4:0] ILA__n19 ; 
    wire[31:0] ILA__n190 ; 
    wire ILA__n191 ; 
    wire[31:0] ILA__n192 ; 
    wire ILA__n193 ; 
    wire[31:0] ILA__n194 ; 
    wire ILA__n195 ; 
    wire[31:0] ILA__n196 ; 
    wire ILA__n197 ; 
    wire[31:0] ILA__n198 ; 
    wire ILA__n199 ; 
    wire ILA__n2 ; 
    wire[31:0] ILA__n200 ; 
    wire ILA__n201 ; 
    wire[31:0] ILA__n202 ; 
    wire ILA__n203 ; 
    wire[31:0] ILA__n204 ; 
    wire ILA__n205 ; 
    wire[31:0] ILA__n206 ; 
    wire ILA__n207 ; 
    wire[31:0] ILA__n208 ; 
    wire ILA__n209 ; 
    wire ILA__n21 ; 
    wire[31:0] ILA__n210 ; 
    wire ILA__n211 ; 
    wire[31:0] ILA__n212 ; 
    wire ILA__n213 ; 
    wire[31:0] ILA__n214 ; 
    wire ILA__n215 ; 
    wire[31:0] ILA__n216 ; 
    wire ILA__n217 ; 
    wire[31:0] ILA__n218 ; 
    wire ILA__n219 ; 
    wire[31:0] ILA__n220 ; 
    wire ILA__n221 ; 
    wire[31:0] ILA__n222 ; 
    wire ILA__n223 ; 
    wire[31:0] ILA__n224 ; 
    wire ILA__n225 ; 
    wire[31:0] ILA__n226 ; 
    wire ILA__n227 ; 
    wire[31:0] ILA__n228 ; 
    wire ILA__n229 ; 
    wire ILA__n23 ; 
    wire[31:0] ILA__n230 ; 
    wire ILA__n231 ; 
    wire[31:0] ILA__n232 ; 
    wire ILA__n233 ; 
    wire[31:0] ILA__n234 ; 
    wire ILA__n235 ; 
    wire[31:0] ILA__n236 ; 
    wire ILA__n25 ; 
    wire ILA__n27 ; 
    wire ILA__n29 ; 
    wire[2:0] ILA__n3 ; 
    wire ILA__n31 ; 
    wire ILA__n33 ; 
    wire ILA__n35 ; 
    wire ILA__n37 ; 
    wire ILA__n39 ; 
    wire ILA__n41 ; 
    wire ILA__n43 ; 
    wire ILA__n45 ; 
    wire ILA__n47 ; 
    wire ILA__n49 ; 
    wire ILA__n5 ; 
    wire ILA__n51 ; 
    wire ILA__n53 ; 
    wire ILA__n55 ; 
    wire ILA__n57 ; 
    wire ILA__n59 ; 
    wire ILA__n6 ; 
    wire ILA__n61 ; 
    wire ILA__n63 ; 
    wire ILA__n65 ; 
    wire ILA__n67 ; 
    wire ILA__n69 ; 
    wire[6:0] ILA__n7 ; 
    wire ILA__n71 ; 
    wire ILA__n73 ; 
    wire ILA__n75 ; 
    wire ILA__n77 ; 
    wire ILA__n79 ; 
    wire ILA__n80 ; 
    wire[31:0] ILA__n81 ; 
    wire[31:0] ILA__n82 ; 
    wire[31:0] ILA__n83 ; 
    wire[31:0] ILA__n84 ; 
    wire[31:0] ILA__n85 ; 
    wire[31:0] ILA__n86 ; 
    wire[31:0] ILA__n87 ; 
    wire[31:0] ILA__n88 ; 
    wire[31:0] ILA__n89 ; 
    wire ILA__n9 ; 
    wire[31:0] ILA__n90 ; 
    wire[31:0] ILA__n91 ; 
    wire[31:0] ILA__n92 ; 
    wire[31:0] ILA__n93 ; 
    wire[31:0] ILA__n94 ; 
    wire[31:0] ILA__n95 ; 
    wire[31:0] ILA__n96 ; 
    wire[31:0] ILA__n97 ; 
    wire[31:0] ILA__n98 ; 
    wire[31:0] ILA__n99 ; (* ILA__keep *)
    wire[31:0] ILA__pc_randinit ; 
    wire ILA__rst ; (* ILA__keep *)
    wire[31:0] ILA__store_addr_randinit ; (* ILA__keep *)
    wire[31:0] ILA__store_data_randinit ; (* ILA__keep *)
    wire ILA__store_en_randinit ; (* ILA__keep *)
    wire[2:0] ILA__store_size_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x0_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x10_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x11_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x12_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x13_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x14_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x15_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x16_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x17_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x18_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x19_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x1_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x20_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x21_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x22_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x23_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x24_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x25_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x26_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x27_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x28_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x29_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x2_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x30_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x31_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x3_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x4_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x5_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x6_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x7_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x8_randinit ; (* ILA__keep *)
    wire[31:0] ILA__x9_randinit ; 
  assign  ILA____ILA_riscv_valid__ =1'b1; 
  assign  ILA__n0 = ILA__inst [6:0]; 
  assign  ILA__bv_7_51_n1 =7'h33; 
  assign  ILA__n2 =( ILA__n0 )==( ILA__bv_7_51_n1 ); 
  assign  ILA__n3 = ILA__inst [14:12]; 
  assign  ILA__bv_3_0_n4 =3'h0; 
  assign  ILA__n5 =( ILA__n3 )==( ILA__bv_3_0_n4 ); 
  assign  ILA__n6 =( ILA__n2 )&( ILA__n5 ); 
  assign  ILA__n7 = ILA__inst [31:25]; 
  assign  ILA__bv_7_0_n8 =7'h0; 
  assign  ILA__n9 =( ILA__n7 )==( ILA__bv_7_0_n8 ); 
  assign  ILA__n10 =( ILA__n6 )&( ILA__n9 ); 
  assign  ILA____ILA_riscv_decode_of_ADD__ = ILA__n10 ; 
  assign  ILA__bv_32_4_n12 =32'h4; 
  assign  ILA__n13 =( ILA__pc )+( ILA__bv_32_4_n12 ); 
  assign  ILA__bv_1_0_n14 =1'h0; 
  assign  ILA__bv_32_0_n15 =32'h0; 
  assign  ILA__n16 = ILA__inst [11:7]; 
  assign  ILA__bv_5_1_n17 =5'h1; 
  assign  ILA__n18 =( ILA__n16 )==( ILA__bv_5_1_n17 ); 
  assign  ILA__n19 = ILA__inst [19:15]; 
  assign  ILA__bv_5_31_n20 =5'h1f; 
  assign  ILA__n21 =( ILA__n19 )==( ILA__bv_5_31_n20 ); 
  assign  ILA__bv_5_30_n22 =5'h1e; 
  assign  ILA__n23 =( ILA__n19 )==( ILA__bv_5_30_n22 ); 
  assign  ILA__bv_5_29_n24 =5'h1d; 
  assign  ILA__n25 =( ILA__n19 )==( ILA__bv_5_29_n24 ); 
  assign  ILA__bv_5_28_n26 =5'h1c; 
  assign  ILA__n27 =( ILA__n19 )==( ILA__bv_5_28_n26 ); 
  assign  ILA__bv_5_27_n28 =5'h1b; 
  assign  ILA__n29 =( ILA__n19 )==( ILA__bv_5_27_n28 ); 
  assign  ILA__bv_5_26_n30 =5'h1a; 
  assign  ILA__n31 =( ILA__n19 )==( ILA__bv_5_26_n30 ); 
  assign  ILA__bv_5_25_n32 =5'h19; 
  assign  ILA__n33 =( ILA__n19 )==( ILA__bv_5_25_n32 ); 
  assign  ILA__bv_5_24_n34 =5'h18; 
  assign  ILA__n35 =( ILA__n19 )==( ILA__bv_5_24_n34 ); 
  assign  ILA__bv_5_23_n36 =5'h17; 
  assign  ILA__n37 =( ILA__n19 )==( ILA__bv_5_23_n36 ); 
  assign  ILA__bv_5_22_n38 =5'h16; 
  assign  ILA__n39 =( ILA__n19 )==( ILA__bv_5_22_n38 ); 
  assign  ILA__bv_5_21_n40 =5'h15; 
  assign  ILA__n41 =( ILA__n19 )==( ILA__bv_5_21_n40 ); 
  assign  ILA__bv_5_20_n42 =5'h14; 
  assign  ILA__n43 =( ILA__n19 )==( ILA__bv_5_20_n42 ); 
  assign  ILA__bv_5_19_n44 =5'h13; 
  assign  ILA__n45 =( ILA__n19 )==( ILA__bv_5_19_n44 ); 
  assign  ILA__bv_5_18_n46 =5'h12; 
  assign  ILA__n47 =( ILA__n19 )==( ILA__bv_5_18_n46 ); 
  assign  ILA__bv_5_17_n48 =5'h11; 
  assign  ILA__n49 =( ILA__n19 )==( ILA__bv_5_17_n48 ); 
  assign  ILA__bv_5_16_n50 =5'h10; 
  assign  ILA__n51 =( ILA__n19 )==( ILA__bv_5_16_n50 ); 
  assign  ILA__bv_5_15_n52 =5'hf; 
  assign  ILA__n53 =( ILA__n19 )==( ILA__bv_5_15_n52 ); 
  assign  ILA__bv_5_14_n54 =5'he; 
  assign  ILA__n55 =( ILA__n19 )==( ILA__bv_5_14_n54 ); 
  assign  ILA__bv_5_13_n56 =5'hd; 
  assign  ILA__n57 =( ILA__n19 )==( ILA__bv_5_13_n56 ); 
  assign  ILA__bv_5_12_n58 =5'hc; 
  assign  ILA__n59 =( ILA__n19 )==( ILA__bv_5_12_n58 ); 
  assign  ILA__bv_5_11_n60 =5'hb; 
  assign  ILA__n61 =( ILA__n19 )==( ILA__bv_5_11_n60 ); 
  assign  ILA__bv_5_10_n62 =5'ha; 
  assign  ILA__n63 =( ILA__n19 )==( ILA__bv_5_10_n62 ); 
  assign  ILA__bv_5_9_n64 =5'h9; 
  assign  ILA__n65 =( ILA__n19 )==( ILA__bv_5_9_n64 ); 
  assign  ILA__bv_5_8_n66 =5'h8; 
  assign  ILA__n67 =( ILA__n19 )==( ILA__bv_5_8_n66 ); 
  assign  ILA__bv_5_7_n68 =5'h7; 
  assign  ILA__n69 =( ILA__n19 )==( ILA__bv_5_7_n68 ); 
  assign  ILA__bv_5_6_n70 =5'h6; 
  assign  ILA__n71 =( ILA__n19 )==( ILA__bv_5_6_n70 ); 
  assign  ILA__bv_5_5_n72 =5'h5; 
  assign  ILA__n73 =( ILA__n19 )==( ILA__bv_5_5_n72 ); 
  assign  ILA__bv_5_4_n74 =5'h4; 
  assign  ILA__n75 =( ILA__n19 )==( ILA__bv_5_4_n74 ); 
  assign  ILA__bv_5_3_n76 =5'h3; 
  assign  ILA__n77 =( ILA__n19 )==( ILA__bv_5_3_n76 ); 
  assign  ILA__bv_5_2_n78 =5'h2; 
  assign  ILA__n79 =( ILA__n19 )==( ILA__bv_5_2_n78 ); 
  assign  ILA__n80 =( ILA__n19 )==( ILA__bv_5_1_n17 ); 
  assign  ILA__n81 =( ILA__n80 ) ? ( ILA__x1 ):( ILA__bv_32_0_n15 ); 
  assign  ILA__n82 =( ILA__n79 ) ? ( ILA__x2 ):( ILA__n81 ); 
  assign  ILA__n83 =( ILA__n77 ) ? ( ILA__x3 ):( ILA__n82 ); 
  assign  ILA__n84 =( ILA__n75 ) ? ( ILA__x4 ):( ILA__n83 ); 
  assign  ILA__n85 =( ILA__n73 ) ? ( ILA__x5 ):( ILA__n84 ); 
  assign  ILA__n86 =( ILA__n71 ) ? ( ILA__x6 ):( ILA__n85 ); 
  assign  ILA__n87 =( ILA__n69 ) ? ( ILA__x7 ):( ILA__n86 ); 
  assign  ILA__n88 =( ILA__n67 ) ? ( ILA__x8 ):( ILA__n87 ); 
  assign  ILA__n89 =( ILA__n65 ) ? ( ILA__x9 ):( ILA__n88 ); 
  assign  ILA__n90 =( ILA__n63 ) ? ( ILA__x10 ):( ILA__n89 ); 
  assign  ILA__n91 =( ILA__n61 ) ? ( ILA__x11 ):( ILA__n90 ); 
  assign  ILA__n92 =( ILA__n59 ) ? ( ILA__x12 ):( ILA__n91 ); 
  assign  ILA__n93 =( ILA__n57 ) ? ( ILA__x13 ):( ILA__n92 ); 
  assign  ILA__n94 =( ILA__n55 ) ? ( ILA__x14 ):( ILA__n93 ); 
  assign  ILA__n95 =( ILA__n53 ) ? ( ILA__x15 ):( ILA__n94 ); 
  assign  ILA__n96 =( ILA__n51 ) ? ( ILA__x16 ):( ILA__n95 ); 
  assign  ILA__n97 =( ILA__n49 ) ? ( ILA__x17 ):( ILA__n96 ); 
  assign  ILA__n98 =( ILA__n47 ) ? ( ILA__x18 ):( ILA__n97 ); 
  assign  ILA__n99 =( ILA__n45 ) ? ( ILA__x19 ):( ILA__n98 ); 
  assign  ILA__n100 =( ILA__n43 ) ? ( ILA__x20 ):( ILA__n99 ); 
  assign  ILA__n101 =( ILA__n41 ) ? ( ILA__x21 ):( ILA__n100 ); 
  assign  ILA__n102 =( ILA__n39 ) ? ( ILA__x22 ):( ILA__n101 ); 
  assign  ILA__n103 =( ILA__n37 ) ? ( ILA__x23 ):( ILA__n102 ); 
  assign  ILA__n104 =( ILA__n35 ) ? ( ILA__x24 ):( ILA__n103 ); 
  assign  ILA__n105 =( ILA__n33 ) ? ( ILA__x25 ):( ILA__n104 ); 
  assign  ILA__n106 =( ILA__n31 ) ? ( ILA__x26 ):( ILA__n105 ); 
  assign  ILA__n107 =( ILA__n29 ) ? ( ILA__x27 ):( ILA__n106 ); 
  assign  ILA__n108 =( ILA__n27 ) ? ( ILA__x28 ):( ILA__n107 ); 
  assign  ILA__n109 =( ILA__n25 ) ? ( ILA__x29 ):( ILA__n108 ); 
  assign  ILA__n110 =( ILA__n23 ) ? ( ILA__x30 ):( ILA__n109 ); 
  assign  ILA__n111 =( ILA__n21 ) ? ( ILA__x31 ):( ILA__n110 ); 
  assign  ILA__n112 = ILA__inst [24:20]; 
  assign  ILA__n113 =( ILA__n112 )==( ILA__bv_5_31_n20 ); 
  assign  ILA__n114 =( ILA__n112 )==( ILA__bv_5_30_n22 ); 
  assign  ILA__n115 =( ILA__n112 )==( ILA__bv_5_29_n24 ); 
  assign  ILA__n116 =( ILA__n112 )==( ILA__bv_5_28_n26 ); 
  assign  ILA__n117 =( ILA__n112 )==( ILA__bv_5_27_n28 ); 
  assign  ILA__n118 =( ILA__n112 )==( ILA__bv_5_26_n30 ); 
  assign  ILA__n119 =( ILA__n112 )==( ILA__bv_5_25_n32 ); 
  assign  ILA__n120 =( ILA__n112 )==( ILA__bv_5_24_n34 ); 
  assign  ILA__n121 =( ILA__n112 )==( ILA__bv_5_23_n36 ); 
  assign  ILA__n122 =( ILA__n112 )==( ILA__bv_5_22_n38 ); 
  assign  ILA__n123 =( ILA__n112 )==( ILA__bv_5_21_n40 ); 
  assign  ILA__n124 =( ILA__n112 )==( ILA__bv_5_20_n42 ); 
  assign  ILA__n125 =( ILA__n112 )==( ILA__bv_5_19_n44 ); 
  assign  ILA__n126 =( ILA__n112 )==( ILA__bv_5_18_n46 ); 
  assign  ILA__n127 =( ILA__n112 )==( ILA__bv_5_17_n48 ); 
  assign  ILA__n128 =( ILA__n112 )==( ILA__bv_5_16_n50 ); 
  assign  ILA__n129 =( ILA__n112 )==( ILA__bv_5_15_n52 ); 
  assign  ILA__n130 =( ILA__n112 )==( ILA__bv_5_14_n54 ); 
  assign  ILA__n131 =( ILA__n112 )==( ILA__bv_5_13_n56 ); 
  assign  ILA__n132 =( ILA__n112 )==( ILA__bv_5_12_n58 ); 
  assign  ILA__n133 =( ILA__n112 )==( ILA__bv_5_11_n60 ); 
  assign  ILA__n134 =( ILA__n112 )==( ILA__bv_5_10_n62 ); 
  assign  ILA__n135 =( ILA__n112 )==( ILA__bv_5_9_n64 ); 
  assign  ILA__n136 =( ILA__n112 )==( ILA__bv_5_8_n66 ); 
  assign  ILA__n137 =( ILA__n112 )==( ILA__bv_5_7_n68 ); 
  assign  ILA__n138 =( ILA__n112 )==( ILA__bv_5_6_n70 ); 
  assign  ILA__n139 =( ILA__n112 )==( ILA__bv_5_5_n72 ); 
  assign  ILA__n140 =( ILA__n112 )==( ILA__bv_5_4_n74 ); 
  assign  ILA__n141 =( ILA__n112 )==( ILA__bv_5_3_n76 ); 
  assign  ILA__n142 =( ILA__n112 )==( ILA__bv_5_2_n78 ); 
  assign  ILA__n143 =( ILA__n112 )==( ILA__bv_5_1_n17 ); 
  assign  ILA__n144 =( ILA__n143 ) ? ( ILA__x1 ):( ILA__bv_32_0_n15 ); 
  assign  ILA__n145 =( ILA__n142 ) ? ( ILA__x2 ):( ILA__n144 ); 
  assign  ILA__n146 =( ILA__n141 ) ? ( ILA__x3 ):( ILA__n145 ); 
  assign  ILA__n147 =( ILA__n140 ) ? ( ILA__x4 ):( ILA__n146 ); 
  assign  ILA__n148 =( ILA__n139 ) ? ( ILA__x5 ):( ILA__n147 ); 
  assign  ILA__n149 =( ILA__n138 ) ? ( ILA__x6 ):( ILA__n148 ); 
  assign  ILA__n150 =( ILA__n137 ) ? ( ILA__x7 ):( ILA__n149 ); 
  assign  ILA__n151 =( ILA__n136 ) ? ( ILA__x8 ):( ILA__n150 ); 
  assign  ILA__n152 =( ILA__n135 ) ? ( ILA__x9 ):( ILA__n151 ); 
  assign  ILA__n153 =( ILA__n134 ) ? ( ILA__x10 ):( ILA__n152 ); 
  assign  ILA__n154 =( ILA__n133 ) ? ( ILA__x11 ):( ILA__n153 ); 
  assign  ILA__n155 =( ILA__n132 ) ? ( ILA__x12 ):( ILA__n154 ); 
  assign  ILA__n156 =( ILA__n131 ) ? ( ILA__x13 ):( ILA__n155 ); 
  assign  ILA__n157 =( ILA__n130 ) ? ( ILA__x14 ):( ILA__n156 ); 
  assign  ILA__n158 =( ILA__n129 ) ? ( ILA__x15 ):( ILA__n157 ); 
  assign  ILA__n159 =( ILA__n128 ) ? ( ILA__x16 ):( ILA__n158 ); 
  assign  ILA__n160 =( ILA__n127 ) ? ( ILA__x17 ):( ILA__n159 ); 
  assign  ILA__n161 =( ILA__n126 ) ? ( ILA__x18 ):( ILA__n160 ); 
  assign  ILA__n162 =( ILA__n125 ) ? ( ILA__x19 ):( ILA__n161 ); 
  assign  ILA__n163 =( ILA__n124 ) ? ( ILA__x20 ):( ILA__n162 ); 
  assign  ILA__n164 =( ILA__n123 ) ? ( ILA__x21 ):( ILA__n163 ); 
  assign  ILA__n165 =( ILA__n122 ) ? ( ILA__x22 ):( ILA__n164 ); 
  assign  ILA__n166 =( ILA__n121 ) ? ( ILA__x23 ):( ILA__n165 ); 
  assign  ILA__n167 =( ILA__n120 ) ? ( ILA__x24 ):( ILA__n166 ); 
  assign  ILA__n168 =( ILA__n119 ) ? ( ILA__x25 ):( ILA__n167 ); 
  assign  ILA__n169 =( ILA__n118 ) ? ( ILA__x26 ):( ILA__n168 ); 
  assign  ILA__n170 =( ILA__n117 ) ? ( ILA__x27 ):( ILA__n169 ); 
  assign  ILA__n171 =( ILA__n116 ) ? ( ILA__x28 ):( ILA__n170 ); 
  assign  ILA__n172 =( ILA__n115 ) ? ( ILA__x29 ):( ILA__n171 ); 
  assign  ILA__n173 =( ILA__n114 ) ? ( ILA__x30 ):( ILA__n172 ); 
  assign  ILA__n174 =( ILA__n113 ) ? ( ILA__x31 ):( ILA__n173 ); 
  assign  ILA__n175 =( ILA__n111 )+( ILA__n174 ); 
  assign  ILA__n176 =( ILA__n18 ) ? ( ILA__n175 ):( ILA__x1 ); 
  assign  ILA__n177 =( ILA__n16 )==( ILA__bv_5_2_n78 ); 
  assign  ILA__n178 =( ILA__n177 ) ? ( ILA__n175 ):( ILA__x2 ); 
  assign  ILA__n179 =( ILA__n16 )==( ILA__bv_5_3_n76 ); 
  assign  ILA__n180 =( ILA__n179 ) ? ( ILA__n175 ):( ILA__x3 ); 
  assign  ILA__n181 =( ILA__n16 )==( ILA__bv_5_4_n74 ); 
  assign  ILA__n182 =( ILA__n181 ) ? ( ILA__n175 ):( ILA__x4 ); 
  assign  ILA__n183 =( ILA__n16 )==( ILA__bv_5_5_n72 ); 
  assign  ILA__n184 =( ILA__n183 ) ? ( ILA__n175 ):( ILA__x5 ); 
  assign  ILA__n185 =( ILA__n16 )==( ILA__bv_5_6_n70 ); 
  assign  ILA__n186 =( ILA__n185 ) ? ( ILA__n175 ):( ILA__x6 ); 
  assign  ILA__n187 =( ILA__n16 )==( ILA__bv_5_7_n68 ); 
  assign  ILA__n188 =( ILA__n187 ) ? ( ILA__n175 ):( ILA__x7 ); 
  assign  ILA__n189 =( ILA__n16 )==( ILA__bv_5_8_n66 ); 
  assign  ILA__n190 =( ILA__n189 ) ? ( ILA__n175 ):( ILA__x8 ); 
  assign  ILA__n191 =( ILA__n16 )==( ILA__bv_5_9_n64 ); 
  assign  ILA__n192 =( ILA__n191 ) ? ( ILA__n175 ):( ILA__x9 ); 
  assign  ILA__n193 =( ILA__n16 )==( ILA__bv_5_10_n62 ); 
  assign  ILA__n194 =( ILA__n193 ) ? ( ILA__n175 ):( ILA__x10 ); 
  assign  ILA__n195 =( ILA__n16 )==( ILA__bv_5_11_n60 ); 
  assign  ILA__n196 =( ILA__n195 ) ? ( ILA__n175 ):( ILA__x11 ); 
  assign  ILA__n197 =( ILA__n16 )==( ILA__bv_5_12_n58 ); 
  assign  ILA__n198 =( ILA__n197 ) ? ( ILA__n175 ):( ILA__x12 ); 
  assign  ILA__n199 =( ILA__n16 )==( ILA__bv_5_13_n56 ); 
  assign  ILA__n200 =( ILA__n199 ) ? ( ILA__n175 ):( ILA__x13 ); 
  assign  ILA__n201 =( ILA__n16 )==( ILA__bv_5_14_n54 ); 
  assign  ILA__n202 =( ILA__n201 ) ? ( ILA__n175 ):( ILA__x14 ); 
  assign  ILA__n203 =( ILA__n16 )==( ILA__bv_5_15_n52 ); 
  assign  ILA__n204 =( ILA__n203 ) ? ( ILA__n175 ):( ILA__x15 ); 
  assign  ILA__n205 =( ILA__n16 )==( ILA__bv_5_16_n50 ); 
  assign  ILA__n206 =( ILA__n205 ) ? ( ILA__n175 ):( ILA__x16 ); 
  assign  ILA__n207 =( ILA__n16 )==( ILA__bv_5_17_n48 ); 
  assign  ILA__n208 =( ILA__n207 ) ? ( ILA__n175 ):( ILA__x17 ); 
  assign  ILA__n209 =( ILA__n16 )==( ILA__bv_5_18_n46 ); 
  assign  ILA__n210 =( ILA__n209 ) ? ( ILA__n175 ):( ILA__x18 ); 
  assign  ILA__n211 =( ILA__n16 )==( ILA__bv_5_19_n44 ); 
  assign  ILA__n212 =( ILA__n211 ) ? ( ILA__n175 ):( ILA__x19 ); 
  assign  ILA__n213 =( ILA__n16 )==( ILA__bv_5_20_n42 ); 
  assign  ILA__n214 =( ILA__n213 ) ? ( ILA__n175 ):( ILA__x20 ); 
  assign  ILA__n215 =( ILA__n16 )==( ILA__bv_5_21_n40 ); 
  assign  ILA__n216 =( ILA__n215 ) ? ( ILA__n175 ):( ILA__x21 ); 
  assign  ILA__n217 =( ILA__n16 )==( ILA__bv_5_22_n38 ); 
  assign  ILA__n218 =( ILA__n217 ) ? ( ILA__n175 ):( ILA__x22 ); 
  assign  ILA__n219 =( ILA__n16 )==( ILA__bv_5_23_n36 ); 
  assign  ILA__n220 =( ILA__n219 ) ? ( ILA__n175 ):( ILA__x23 ); 
  assign  ILA__n221 =( ILA__n16 )==( ILA__bv_5_24_n34 ); 
  assign  ILA__n222 =( ILA__n221 ) ? ( ILA__n175 ):( ILA__x24 ); 
  assign  ILA__n223 =( ILA__n16 )==( ILA__bv_5_25_n32 ); 
  assign  ILA__n224 =( ILA__n223 ) ? ( ILA__n175 ):( ILA__x25 ); 
  assign  ILA__n225 =( ILA__n16 )==( ILA__bv_5_26_n30 ); 
  assign  ILA__n226 =( ILA__n225 ) ? ( ILA__n175 ):( ILA__x26 ); 
  assign  ILA__n227 =( ILA__n16 )==( ILA__bv_5_27_n28 ); 
  assign  ILA__n228 =( ILA__n227 ) ? ( ILA__n175 ):( ILA__x27 ); 
  assign  ILA__n229 =( ILA__n16 )==( ILA__bv_5_28_n26 ); 
  assign  ILA__n230 =( ILA__n229 ) ? ( ILA__n175 ):( ILA__x28 ); 
  assign  ILA__n231 =( ILA__n16 )==( ILA__bv_5_29_n24 ); 
  assign  ILA__n232 =( ILA__n231 ) ? ( ILA__n175 ):( ILA__x29 ); 
  assign  ILA__n233 =( ILA__n16 )==( ILA__bv_5_30_n22 ); 
  assign  ILA__n234 =( ILA__n233 ) ? ( ILA__n175 ):( ILA__x30 ); 
  assign  ILA__n235 =( ILA__n16 )==( ILA__bv_5_31_n20 ); 
  assign  ILA__n236 =( ILA__n235 ) ? ( ILA__n175 ):( ILA__x31 ); 
  always @( posedge  ILA__clk )
         begin 
             if ( ILA__rst )
                 begin  
                     ILA__pc  <= ILA__pc_randinit ; 
                     ILA__load_en  <= ILA__load_en_randinit ; 
                     ILA__load_addr  <= ILA__load_addr_randinit ; 
                     ILA__load_size  <= ILA__load_size_randinit ; 
                     ILA__load_data  <= ILA__load_data_randinit ; 
                     ILA__store_en  <= ILA__store_en_randinit ; 
                     ILA__store_addr  <= ILA__store_addr_randinit ; 
                     ILA__store_size  <= ILA__store_size_randinit ; 
                     ILA__store_data  <= ILA__store_data_randinit ; 
                     ILA__x0  <= ILA__x0_randinit ; 
                     ILA__x1  <= ILA__x1_randinit ; 
                     ILA__x2  <= ILA__x2_randinit ; 
                     ILA__x3  <= ILA__x3_randinit ; 
                     ILA__x4  <= ILA__x4_randinit ; 
                     ILA__x5  <= ILA__x5_randinit ; 
                     ILA__x6  <= ILA__x6_randinit ; 
                     ILA__x7  <= ILA__x7_randinit ; 
                     ILA__x8  <= ILA__x8_randinit ; 
                     ILA__x9  <= ILA__x9_randinit ; 
                     ILA__x10  <= ILA__x10_randinit ; 
                     ILA__x11  <= ILA__x11_randinit ; 
                     ILA__x12  <= ILA__x12_randinit ; 
                     ILA__x13  <= ILA__x13_randinit ; 
                     ILA__x14  <= ILA__x14_randinit ; 
                     ILA__x15  <= ILA__x15_randinit ; 
                     ILA__x16  <= ILA__x16_randinit ; 
                     ILA__x17  <= ILA__x17_randinit ; 
                     ILA__x18  <= ILA__x18_randinit ; 
                     ILA__x19  <= ILA__x19_randinit ; 
                     ILA__x20  <= ILA__x20_randinit ; 
                     ILA__x21  <= ILA__x21_randinit ; 
                     ILA__x22  <= ILA__x22_randinit ; 
                     ILA__x23  <= ILA__x23_randinit ; 
                     ILA__x24  <= ILA__x24_randinit ; 
                     ILA__x25  <= ILA__x25_randinit ; 
                     ILA__x26  <= ILA__x26_randinit ; 
                     ILA__x27  <= ILA__x27_randinit ; 
                     ILA__x28  <= ILA__x28_randinit ; 
                     ILA__x29  <= ILA__x29_randinit ; 
                     ILA__x30  <= ILA__x30_randinit ; 
                     ILA__x31  <= ILA__x31_randinit ; 
                     ILA____COUNTER_start__n11  <=0;
                 end 
              else 
                 if ( ILA____START__ && ILA____ILA_riscv_valid__ )
                     begin 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA____COUNTER_start__n11  <=1;
                             end 
                          else 
                             if (( ILA____COUNTER_start__n11 >=1)&&( ILA____COUNTER_start__n11 <255))
                                 begin  
                                     ILA____COUNTER_start__n11  <= ILA____COUNTER_start__n11 +1;
                                 end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__pc  <= ILA__n13 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__load_en  <= ILA__bv_1_0_n14 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__load_addr  <= ILA__load_addr ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__load_size  <= ILA__load_size ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__load_data  <= ILA__load_data ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__store_en  <= ILA__bv_1_0_n14 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__store_addr  <= ILA__store_addr ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__store_size  <= ILA__store_size ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__store_data  <= ILA__store_data ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x0  <= ILA__bv_32_0_n15 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x1  <= ILA__n176 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x2  <= ILA__n178 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x3  <= ILA__n180 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x4  <= ILA__n182 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x5  <= ILA__n184 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x6  <= ILA__n186 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x7  <= ILA__n188 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x8  <= ILA__n190 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x9  <= ILA__n192 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x10  <= ILA__n194 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x11  <= ILA__n196 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x12  <= ILA__n198 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x13  <= ILA__n200 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x14  <= ILA__n202 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x15  <= ILA__n204 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x16  <= ILA__n206 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x17  <= ILA__n208 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x18  <= ILA__n210 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x19  <= ILA__n212 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x20  <= ILA__n214 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x21  <= ILA__n216 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x22  <= ILA__n218 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x23  <= ILA__n220 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x24  <= ILA__n222 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x25  <= ILA__n224 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x26  <= ILA__n226 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x27  <= ILA__n228 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x28  <= ILA__n230 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x29  <= ILA__n232 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x30  <= ILA__n234 ;
                             end 
                         if ( ILA____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA__x31  <= ILA__n236 ;
                             end 
                     end 
         end
 
    assign ILA____START__ = __START__;
    assign ILA__clk = clk;
    assign ILA__inst = __ILA_I_inst;
    assign ILA__rst = rst;
    assign __ILA_riscv_decode_of_ADD__ = ILA____ILA_riscv_decode_of_ADD__;
    assign __ILA_riscv_valid__ = ILA____ILA_riscv_valid__;
    assign __ILA_SO_pc = ILA__pc;
    assign __ILA_SO_load_en = ILA__load_en;
    assign __ILA_SO_load_addr = ILA__load_addr;
    assign __ILA_SO_load_size = ILA__load_size;
    assign __ILA_SO_load_data = ILA__load_data;
    assign __ILA_SO_store_en = ILA__store_en;
    assign __ILA_SO_store_addr = ILA__store_addr;
    assign __ILA_SO_store_size = ILA__store_size;
    assign __ILA_SO_store_data = ILA__store_data;
    assign __ILA_SO_x0 = ILA__x0;
    assign __ILA_SO_x1 = ILA__x1;
    assign __ILA_SO_x2 = ILA__x2;
    assign __ILA_SO_x3 = ILA__x3;
    assign __ILA_SO_x4 = ILA__x4;
    assign __ILA_SO_x5 = ILA__x5;
    assign __ILA_SO_x6 = ILA__x6;
    assign __ILA_SO_x7 = ILA__x7;
    assign __ILA_SO_x8 = ILA__x8;
    assign __ILA_SO_x9 = ILA__x9;
    assign __ILA_SO_x10 = ILA__x10;
    assign __ILA_SO_x11 = ILA__x11;
    assign __ILA_SO_x12 = ILA__x12;
    assign __ILA_SO_x13 = ILA__x13;
    assign __ILA_SO_x14 = ILA__x14;
    assign __ILA_SO_x15 = ILA__x15;
    assign __ILA_SO_x16 = ILA__x16;
    assign __ILA_SO_x17 = ILA__x17;
    assign __ILA_SO_x18 = ILA__x18;
    assign __ILA_SO_x19 = ILA__x19;
    assign __ILA_SO_x20 = ILA__x20;
    assign __ILA_SO_x21 = ILA__x21;
    assign __ILA_SO_x22 = ILA__x22;
    assign __ILA_SO_x23 = ILA__x23;
    assign __ILA_SO_x24 = ILA__x24;
    assign __ILA_SO_x25 = ILA__x25;
    assign __ILA_SO_x26 = ILA__x26;
    assign __ILA_SO_x27 = ILA__x27;
    assign __ILA_SO_x28 = ILA__x28;
    assign __ILA_SO_x29 = ILA__x29;
    assign __ILA_SO_x30 = ILA__x30;
    assign __ILA_SO_x31 = ILA__x31;
    
assign __EDCOND__ = (end_of_pipeline)&&(__STARTED__) ;
assign __IEND__ = ((((end_of_pipeline)&&(__STARTED__))&&(__RESETED__))&&(!(__ENDED__)))&&(1'b1) ;
assign __VLG_II_m_external_interrupt_req_set_not_clear = 1'b0 ;
assign __VLG_II_nmi_req_set_not_clear = 1'b0 ;
assign __VLG_II_s_external_interrupt_req_set_not_clear = 1'b0 ;
assign __VLG_II_software_interrupt_req_set_not_clear = 1'b0 ;
assign __VLG_II_timer_interrupt_req_set_not_clear = 1'b0 ;
assign __auxvar10__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar10__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ ;
assign __auxvar11__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar11__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ ;
assign __auxvar12__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar12__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ ;
assign __auxvar13__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar13__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ ;
assign __auxvar14__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar14__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ ;
assign __auxvar15__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar15__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ ;
assign __auxvar16__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar16__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ ;
assign __auxvar17__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar17__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ ;
assign __auxvar18__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar18__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ ;
assign __auxvar19__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar19__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ ;
assign __auxvar1__recorder_sn_cond = ((monitor_s2)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar1__recorder_sn_value = RTL__DOT__near_mem$imem_pc ;
assign __auxvar20__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar20__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ ;
assign __auxvar21__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar21__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ ;
assign __auxvar22__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar22__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ ;
assign __auxvar23__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar23__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ ;
assign __auxvar24__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar24__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ ;
assign __auxvar25__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar25__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ ;
assign __auxvar26__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar26__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ ;
assign __auxvar27__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar27__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ ;
assign __auxvar28__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar28__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ ;
assign __auxvar29__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar29__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ ;
assign __auxvar2__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar2__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ ;
assign __auxvar30__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar30__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ ;
assign __auxvar31__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar31__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ ;
assign __auxvar32__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar32__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ ;
assign __auxvar33__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar33__recorder_sn_value = RTL__DOT__near_mem$dmem_req_addr ;
assign __auxvar34__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar34__recorder_sn_value = RTL__DOT__near_mem$EN_dmem_req ;
assign __auxvar35__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar35__recorder_sn_value = RTL__DOT__near_mem$dmem_req_f3 ;
assign __auxvar36__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar36__recorder_sn_value = RTL__DOT__near_mem$dmem_req_op ;
assign __auxvar37__recorder_sn_cond = ((monitor_s2)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar37__recorder_sn_value = RTL__DOT__near_mem$dmem_word64[31:0] ;
assign __auxvar38__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar38__recorder_sn_value = RTL__DOT__near_mem$dmem_req_store_value[31:0] ;
assign __auxvar3__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar3__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ ;
assign __auxvar4__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar4__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ ;
assign __auxvar5__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar5__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ ;
assign __auxvar6__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar6__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ ;
assign __auxvar7__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar7__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ ;
assign __auxvar8__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar8__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ ;
assign __auxvar9__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar9__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ ;
assign __auxvar0__delay_d_0 = monitor_s4 ;
assign end_of_pipeline = (monitor_s4)&&(~(__auxvar0__delay)) ;
assign monitor_s1 = ((RTL__DOT__stage1_rg_full)&(~(monitor_s1_already)))&(__START__) ;
assign s2_enter = ((RTL__DOT__s1_to_s2$D_IN)&(RTL__DOT__s1_to_s2$EN))&(monitor_s1) ;
assign s2_exit = (RTL__DOT__s2_to_s3$D_IN)&(RTL__DOT__s2_to_s3$EN) ;
assign s3_enter = ((RTL__DOT__s2_to_s3$D_IN)&(RTL__DOT__s2_to_s3$EN))&(monitor_s2) ;
assign s3_exit = (RTL__DOT__s3_deq$EN)&(RTL__DOT__s3_deq$D_IN) ;
assign s4_enter = (monitor_s3)&&(RTL__DOT__rg_retiring$EN) ;
assign monitor_s1_already_enter_cond = (monitor_s1)&&(s2_enter) ;
assign monitor_s2_enter_cond = s2_enter ;
assign monitor_s2_exit_cond = s2_exit ;
assign monitor_s3_enter_cond = s3_enter ;
assign monitor_s3_exit_cond = s3_exit ;
assign monitor_s4_enter_cond = s4_enter ;
assign mem_req_addr = __auxvar33__recorder ;
assign mem_req_en = __auxvar34__recorder ;
assign mem_req_funct3 = __auxvar35__recorder ;
assign mem_req_op = __auxvar36__recorder ;
assign mem_req_rd_data = __auxvar37__recorder ;
assign mem_req_wd_data = __auxvar38__recorder ;
assign input_map_assume___p0__ = (!(__START__))||((__ILA_I_inst)==(RTL__DOT__near_mem$imem_instr)) ;
assign invariant_assume__p1__ = !(((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p2__ = !(((RTL__DOT__f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p3__ = !(((RTL__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p4__ = !(((RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p5__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p6__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p7__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p8__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg)==(0))) ;
assign invariant_assume__p9__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p10__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg)==(0))) ;
assign invariant_assume__p11__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p12__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg)==(0))) ;
assign invariant_assume__p13__ = !(((RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p14__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p15__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p16__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p17__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg)==(0))) ;
assign invariant_assume__p18__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p19__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg)==(0))) ;
assign invariant_assume__p20__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p21__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg)==(0))) ;
assign invariant_assume__p22__ = !(((RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__stage1_f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p23__ = !(((RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__stage1_f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p24__ = !(((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__stage2_f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p25__ = !(((RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__stage2_f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p26__ = !(((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p27__ = !(((RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p28__ = ((((!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1)))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__stage3_rg_full)==(1'b1))))&&((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__f_reset_reqs__DOT__full_reg)==(1'b0)))))&&(((!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1)))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__stage2_rg_full)==(1'b1)))) ;
assign invariant_assume__p29__ = ((!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1))))&&((RTL__DOT__stage2_f_reset_reqs__DOT__full_reg)==(1'b1)) ;
assign invariant_assume__p30__ = (((!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1)))||(!((RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg)==(1'b0))))||(!((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(1'b0))))&&((((!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1)))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg)==(1'b0)))) ;
assign invariant_assume__p31__ = (((((((((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b1))))||(!((RTL__DOT__rg_run_on_reset)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!(RTL__DOT__stage2_rg_stage2[101:101])))||((RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr[4:4])==(1'b1)))||(!((RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa[4:4])==(1'b1))))&&(!((RTL__DOT__csr_regfile__DOT__rg_nmi)==(1'b1))))&&(((!((RTL__DOT__rg_state[0:0])==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b0)))))&&(((((((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(1'b1))||(!(RTL__DOT__rg_trap_instr[22:22])))||(!(RTL__DOT__rg_trap_instr[20:20])))||(!(RTL__DOT__rg_trap_instr[26:26])))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b0)))))&&(((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__rg_run_on_reset)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(1'b0)))) ;
assign invariant_assume__p32__ = (((((!((RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg)==(1'b0)))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(1'b0))))&&(((((!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0)))||(!((RTL__DOT__rg_state[0:0])==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(RTL__DOT__rg_run_on_reset)))&&(((((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__rg_state[0:0])==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(RTL__DOT__stage2_rg_stage2[168:168]))||(!(RTL__DOT__rg_cur_priv[1:1]))) ;
assign issue_decode__p33__ = (!(__START__))||(__ILA_riscv_decode_of_ADD__) ;
assign issue_valid__p34__ = (!(__START__))||(__ILA_riscv_valid__) ;
assign noreset__p35__ = (!(__RESETED__))||(!(dummy_reset)) ;
assign post_value_holder__p36__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar10__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar10__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_)) ;
assign post_value_holder__p37__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar11__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar11__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_)) ;
assign post_value_holder__p38__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar12__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar12__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_)) ;
assign post_value_holder__p39__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar13__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar13__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_)) ;
assign post_value_holder__p40__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar14__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar14__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_)) ;
assign post_value_holder__p41__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar15__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar15__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_)) ;
assign post_value_holder__p42__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar16__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar16__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_)) ;
assign post_value_holder__p43__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar17__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar17__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_)) ;
assign post_value_holder__p44__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar18__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar18__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_)) ;
assign post_value_holder__p45__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar19__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar19__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_)) ;
assign post_value_holder__p46__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar1__recorder_sn_condmet)))&&(monitor_s2)))||((__auxvar1__recorder)==(RTL__DOT__near_mem$imem_pc)) ;
assign post_value_holder__p47__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar20__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar20__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_)) ;
assign post_value_holder__p48__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar21__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar21__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_)) ;
assign post_value_holder__p49__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar22__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar22__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_)) ;
assign post_value_holder__p50__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar23__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar23__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_)) ;
assign post_value_holder__p51__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar24__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar24__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_)) ;
assign post_value_holder__p52__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar25__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar25__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_)) ;
assign post_value_holder__p53__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar26__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar26__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_)) ;
assign post_value_holder__p54__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar27__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar27__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_)) ;
assign post_value_holder__p55__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar28__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar28__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_)) ;
assign post_value_holder__p56__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar29__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar29__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_)) ;
assign post_value_holder__p57__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar2__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar2__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_)) ;
assign post_value_holder__p58__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar30__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar30__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_)) ;
assign post_value_holder__p59__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar31__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar31__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_)) ;
assign post_value_holder__p60__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar32__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar32__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_)) ;
assign post_value_holder__p61__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar33__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar33__recorder)==(RTL__DOT__near_mem$dmem_req_addr)) ;
assign post_value_holder__p62__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar34__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar34__recorder)==(RTL__DOT__near_mem$EN_dmem_req)) ;
assign post_value_holder__p63__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar35__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar35__recorder)==(RTL__DOT__near_mem$dmem_req_f3)) ;
assign post_value_holder__p64__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar36__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar36__recorder)==(RTL__DOT__near_mem$dmem_req_op)) ;
assign post_value_holder__p65__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar37__recorder_sn_condmet)))&&(monitor_s2)))||((__auxvar37__recorder)==(RTL__DOT__near_mem$dmem_word64[31:0])) ;
assign post_value_holder__p66__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar38__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar38__recorder)==(RTL__DOT__near_mem$dmem_req_store_value[31:0])) ;
assign post_value_holder__p67__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar3__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar3__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_)) ;
assign post_value_holder__p68__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar4__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar4__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_)) ;
assign post_value_holder__p69__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar5__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar5__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_)) ;
assign post_value_holder__p70__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar6__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar6__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_)) ;
assign post_value_holder__p71__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar7__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar7__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_)) ;
assign post_value_holder__p72__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar8__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar8__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_)) ;
assign post_value_holder__p73__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar9__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar9__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_)) ;
assign rfassumptions__p74__ = (__ILA_SO_pc[1:0])==(2'b00) ;
assign rfassumptions__p75__ = (RTL__DOT__near_mem$imem_pc[1:0])==(2'b00) ;
assign rfassumptions__p76__ = (!(monitor_s2))||((RTL__DOT__near_mem$dmem_exc)==(0)) ;
assign variable_map_assume___p77__ = (!(__START__))||((!((__IEND__)&&(__ILA_SO_load_en)))||((__ILA_SO_load_addr)==(mem_req_addr))) ;
assign variable_map_assume___p78__ = (!(__START__))||((!((__START__)&&(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b0)))))||((__ILA_SO_load_data)==(mem_req_rd_data))) ;
assign variable_map_assume___p79__ = (!(__START__))||((!(__IEND__))||((__ILA_SO_load_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b0))))) ;
assign variable_map_assume___p80__ = (!(__START__))||(((((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))||(((mem_req_funct3)==(0))||((mem_req_funct3)==(4))))&&((!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2)))))||(((mem_req_funct3)==(1))||((mem_req_funct3)==(5)))))&&((!(((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(4)))))||(((mem_req_funct3)==(2))||((mem_req_funct3)==(6)))))&&((!((((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2))))))&&(!(((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(4))))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(8)))))||((mem_req_funct3)==(3)))) ;
assign variable_map_assume___p81__ = (!(__START__))||(((!(__START__))||((__ILA_SO_pc)==(RTL__DOT__near_mem$imem_pc)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_pc)==(__auxvar1__recorder)))) ;
assign variable_map_assume___p82__ = (!(__START__))||((!((__IEND__)&&(__ILA_SO_store_en)))||((__ILA_SO_store_addr)==(mem_req_addr))) ;
assign variable_map_assume___p83__ = (!(__START__))||((!((__IEND__)&&(__ILA_SO_store_en)))||((__ILA_SO_store_data)==(mem_req_wd_data))) ;
assign variable_map_assume___p84__ = (!(__START__))||((!(__IEND__))||((__ILA_SO_store_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b1))))) ;
assign variable_map_assume___p85__ = (!(__START__))||(((((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))||(((mem_req_funct3)==(0))||((mem_req_funct3)==(4))))&&((!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2)))))||(((mem_req_funct3)==(1))||((mem_req_funct3)==(5)))))&&((!(((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(4)))))||(((mem_req_funct3)==(2))||((mem_req_funct3)==(6)))))&&((!((((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2))))))&&(!(((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(4))))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(8)))))||((mem_req_funct3)==(3)))) ;
assign variable_map_assume___p86__ = (!(__START__))||((__ILA_SO_x0)==(0)) ;
assign variable_map_assume___p87__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x1)==(__auxvar2__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x1)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_)))) ;
assign variable_map_assume___p88__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x10)==(__auxvar3__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x10)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_)))) ;
assign variable_map_assume___p89__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x11)==(__auxvar4__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x11)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_)))) ;
assign variable_map_assume___p90__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x12)==(__auxvar5__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x12)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_)))) ;
assign variable_map_assume___p91__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x13)==(__auxvar6__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x13)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_)))) ;
assign variable_map_assume___p92__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x14)==(__auxvar7__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x14)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_)))) ;
assign variable_map_assume___p93__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x15)==(__auxvar8__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x15)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_)))) ;
assign variable_map_assume___p94__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x16)==(__auxvar9__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x16)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_)))) ;
assign variable_map_assume___p95__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x17)==(__auxvar10__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x17)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_)))) ;
assign variable_map_assume___p96__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x18)==(__auxvar11__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x18)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_)))) ;
assign variable_map_assume___p97__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x19)==(__auxvar12__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x19)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_)))) ;
assign variable_map_assume___p98__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x2)==(__auxvar13__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x2)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_)))) ;
assign variable_map_assume___p99__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x20)==(__auxvar14__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x20)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_)))) ;
assign variable_map_assume___p100__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x21)==(__auxvar15__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x21)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_)))) ;
assign variable_map_assume___p101__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x22)==(__auxvar16__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x22)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_)))) ;
assign variable_map_assume___p102__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x23)==(__auxvar17__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x23)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_)))) ;
assign variable_map_assume___p103__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x24)==(__auxvar18__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x24)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_)))) ;
assign variable_map_assume___p104__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x25)==(__auxvar19__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x25)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_)))) ;
assign variable_map_assume___p105__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x26)==(__auxvar20__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x26)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_)))) ;
assign variable_map_assume___p106__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x27)==(__auxvar21__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x27)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_)))) ;
assign variable_map_assume___p107__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x28)==(__auxvar22__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x28)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_)))) ;
assign variable_map_assume___p108__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x29)==(__auxvar23__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x29)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_)))) ;
assign variable_map_assume___p109__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x3)==(__auxvar24__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x3)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_)))) ;
assign variable_map_assume___p110__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x30)==(__auxvar25__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x30)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_)))) ;
assign variable_map_assume___p111__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x31)==(__auxvar26__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x31)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_)))) ;
assign variable_map_assume___p112__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x4)==(__auxvar27__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x4)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_)))) ;
assign variable_map_assume___p113__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x5)==(__auxvar28__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x5)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_)))) ;
assign variable_map_assume___p114__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x6)==(__auxvar29__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x6)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_)))) ;
assign variable_map_assume___p115__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x7)==(__auxvar30__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x7)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_)))) ;
assign variable_map_assume___p116__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x8)==(__auxvar31__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x8)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_)))) ;
assign variable_map_assume___p117__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x9)==(__auxvar32__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x9)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_)))) ;
assign variable_map_assert__p118__ = (!(__IEND__))||((!(__IEND__))||((__ILA_SO_load_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b0))))) ;
assign variable_map_assert__p119__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_pc)==(RTL__DOT__near_mem$imem_pc)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_pc)==(__auxvar1__recorder)))) ;
assign variable_map_assert__p120__ = (!(__IEND__))||((!(__IEND__))||((__ILA_SO_store_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b1))))) ;
assign variable_map_assert__p121__ = (!(__IEND__))||((__ILA_SO_x0)==(0)) ;
assign variable_map_assert__p122__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x1)==(__auxvar2__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x1)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_)))) ;
assign variable_map_assert__p123__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x10)==(__auxvar3__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x10)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_)))) ;
assign variable_map_assert__p124__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x11)==(__auxvar4__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x11)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_)))) ;
assign variable_map_assert__p125__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x12)==(__auxvar5__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x12)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_)))) ;
assign variable_map_assert__p126__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x13)==(__auxvar6__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x13)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_)))) ;
assign variable_map_assert__p127__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x14)==(__auxvar7__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x14)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_)))) ;
assign variable_map_assert__p128__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x15)==(__auxvar8__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x15)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_)))) ;
assign variable_map_assert__p129__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x16)==(__auxvar9__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x16)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_)))) ;
assign variable_map_assert__p130__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x17)==(__auxvar10__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x17)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_)))) ;
assign variable_map_assert__p131__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x18)==(__auxvar11__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x18)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_)))) ;
assign variable_map_assert__p132__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x19)==(__auxvar12__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x19)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_)))) ;
assign variable_map_assert__p133__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x2)==(__auxvar13__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x2)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_)))) ;
assign variable_map_assert__p134__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x20)==(__auxvar14__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x20)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_)))) ;
assign variable_map_assert__p135__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x21)==(__auxvar15__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x21)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_)))) ;
assign variable_map_assert__p136__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x22)==(__auxvar16__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x22)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_)))) ;
assign variable_map_assert__p137__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x23)==(__auxvar17__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x23)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_)))) ;
assign variable_map_assert__p138__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x24)==(__auxvar18__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x24)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_)))) ;
assign variable_map_assert__p139__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x25)==(__auxvar19__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x25)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_)))) ;
assign variable_map_assert__p140__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x26)==(__auxvar20__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x26)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_)))) ;
assign variable_map_assert__p141__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x27)==(__auxvar21__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x27)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_)))) ;
assign variable_map_assert__p142__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x28)==(__auxvar22__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x28)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_)))) ;
assign variable_map_assert__p143__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x29)==(__auxvar23__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x29)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_)))) ;
assign variable_map_assert__p144__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x3)==(__auxvar24__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x3)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_)))) ;
assign variable_map_assert__p145__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x30)==(__auxvar25__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x30)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_)))) ;
assign variable_map_assert__p146__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x31)==(__auxvar26__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x31)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_)))) ;
assign variable_map_assert__p147__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x4)==(__auxvar27__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x4)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_)))) ;
assign variable_map_assert__p148__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x5)==(__auxvar28__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x5)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_)))) ;
assign variable_map_assert__p149__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x6)==(__auxvar29__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x6)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_)))) ;
assign variable_map_assert__p150__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x7)==(__auxvar30__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x7)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_)))) ;
assign variable_map_assert__p151__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x8)==(__auxvar31__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x8)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_)))) ;
assign variable_map_assert__p152__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x9)==(__auxvar32__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x9)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_)))) ;
assign post_value_holder_overly_constrained__p153__ = (!((__auxvar10__recorder_sn_condmet)&&(__auxvar10__recorder_sn_cond)))||((__auxvar10__recorder_sn_value)==(__auxvar10__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p154__ = (!((__auxvar11__recorder_sn_condmet)&&(__auxvar11__recorder_sn_cond)))||((__auxvar11__recorder_sn_value)==(__auxvar11__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p155__ = (!((__auxvar12__recorder_sn_condmet)&&(__auxvar12__recorder_sn_cond)))||((__auxvar12__recorder_sn_value)==(__auxvar12__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p156__ = (!((__auxvar13__recorder_sn_condmet)&&(__auxvar13__recorder_sn_cond)))||((__auxvar13__recorder_sn_value)==(__auxvar13__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p157__ = (!((__auxvar14__recorder_sn_condmet)&&(__auxvar14__recorder_sn_cond)))||((__auxvar14__recorder_sn_value)==(__auxvar14__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p158__ = (!((__auxvar15__recorder_sn_condmet)&&(__auxvar15__recorder_sn_cond)))||((__auxvar15__recorder_sn_value)==(__auxvar15__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p159__ = (!((__auxvar16__recorder_sn_condmet)&&(__auxvar16__recorder_sn_cond)))||((__auxvar16__recorder_sn_value)==(__auxvar16__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p160__ = (!((__auxvar17__recorder_sn_condmet)&&(__auxvar17__recorder_sn_cond)))||((__auxvar17__recorder_sn_value)==(__auxvar17__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p161__ = (!((__auxvar18__recorder_sn_condmet)&&(__auxvar18__recorder_sn_cond)))||((__auxvar18__recorder_sn_value)==(__auxvar18__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p162__ = (!((__auxvar19__recorder_sn_condmet)&&(__auxvar19__recorder_sn_cond)))||((__auxvar19__recorder_sn_value)==(__auxvar19__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p163__ = (!((__auxvar1__recorder_sn_condmet)&&(__auxvar1__recorder_sn_cond)))||((__auxvar1__recorder_sn_value)==(__auxvar1__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p164__ = (!((__auxvar20__recorder_sn_condmet)&&(__auxvar20__recorder_sn_cond)))||((__auxvar20__recorder_sn_value)==(__auxvar20__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p165__ = (!((__auxvar21__recorder_sn_condmet)&&(__auxvar21__recorder_sn_cond)))||((__auxvar21__recorder_sn_value)==(__auxvar21__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p166__ = (!((__auxvar22__recorder_sn_condmet)&&(__auxvar22__recorder_sn_cond)))||((__auxvar22__recorder_sn_value)==(__auxvar22__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p167__ = (!((__auxvar23__recorder_sn_condmet)&&(__auxvar23__recorder_sn_cond)))||((__auxvar23__recorder_sn_value)==(__auxvar23__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p168__ = (!((__auxvar24__recorder_sn_condmet)&&(__auxvar24__recorder_sn_cond)))||((__auxvar24__recorder_sn_value)==(__auxvar24__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p169__ = (!((__auxvar25__recorder_sn_condmet)&&(__auxvar25__recorder_sn_cond)))||((__auxvar25__recorder_sn_value)==(__auxvar25__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p170__ = (!((__auxvar26__recorder_sn_condmet)&&(__auxvar26__recorder_sn_cond)))||((__auxvar26__recorder_sn_value)==(__auxvar26__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p171__ = (!((__auxvar27__recorder_sn_condmet)&&(__auxvar27__recorder_sn_cond)))||((__auxvar27__recorder_sn_value)==(__auxvar27__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p172__ = (!((__auxvar28__recorder_sn_condmet)&&(__auxvar28__recorder_sn_cond)))||((__auxvar28__recorder_sn_value)==(__auxvar28__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p173__ = (!((__auxvar29__recorder_sn_condmet)&&(__auxvar29__recorder_sn_cond)))||((__auxvar29__recorder_sn_value)==(__auxvar29__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p174__ = (!((__auxvar2__recorder_sn_condmet)&&(__auxvar2__recorder_sn_cond)))||((__auxvar2__recorder_sn_value)==(__auxvar2__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p175__ = (!((__auxvar30__recorder_sn_condmet)&&(__auxvar30__recorder_sn_cond)))||((__auxvar30__recorder_sn_value)==(__auxvar30__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p176__ = (!((__auxvar31__recorder_sn_condmet)&&(__auxvar31__recorder_sn_cond)))||((__auxvar31__recorder_sn_value)==(__auxvar31__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p177__ = (!((__auxvar32__recorder_sn_condmet)&&(__auxvar32__recorder_sn_cond)))||((__auxvar32__recorder_sn_value)==(__auxvar32__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p178__ = (!((__auxvar33__recorder_sn_condmet)&&(__auxvar33__recorder_sn_cond)))||((__auxvar33__recorder_sn_value)==(__auxvar33__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p179__ = (!((__auxvar34__recorder_sn_condmet)&&(__auxvar34__recorder_sn_cond)))||((__auxvar34__recorder_sn_value)==(__auxvar34__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p180__ = (!((__auxvar35__recorder_sn_condmet)&&(__auxvar35__recorder_sn_cond)))||((__auxvar35__recorder_sn_value)==(__auxvar35__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p181__ = (!((__auxvar36__recorder_sn_condmet)&&(__auxvar36__recorder_sn_cond)))||((__auxvar36__recorder_sn_value)==(__auxvar36__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p182__ = (!((__auxvar37__recorder_sn_condmet)&&(__auxvar37__recorder_sn_cond)))||((__auxvar37__recorder_sn_value)==(__auxvar37__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p183__ = (!((__auxvar38__recorder_sn_condmet)&&(__auxvar38__recorder_sn_cond)))||((__auxvar38__recorder_sn_value)==(__auxvar38__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p184__ = (!((__auxvar3__recorder_sn_condmet)&&(__auxvar3__recorder_sn_cond)))||((__auxvar3__recorder_sn_value)==(__auxvar3__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p185__ = (!((__auxvar4__recorder_sn_condmet)&&(__auxvar4__recorder_sn_cond)))||((__auxvar4__recorder_sn_value)==(__auxvar4__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p186__ = (!((__auxvar5__recorder_sn_condmet)&&(__auxvar5__recorder_sn_cond)))||((__auxvar5__recorder_sn_value)==(__auxvar5__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p187__ = (!((__auxvar6__recorder_sn_condmet)&&(__auxvar6__recorder_sn_cond)))||((__auxvar6__recorder_sn_value)==(__auxvar6__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p188__ = (!((__auxvar7__recorder_sn_condmet)&&(__auxvar7__recorder_sn_cond)))||((__auxvar7__recorder_sn_value)==(__auxvar7__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p189__ = (!((__auxvar8__recorder_sn_condmet)&&(__auxvar8__recorder_sn_cond)))||((__auxvar8__recorder_sn_value)==(__auxvar8__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p190__ = (!((__auxvar9__recorder_sn_condmet)&&(__auxvar9__recorder_sn_cond)))||((__auxvar9__recorder_sn_value)==(__auxvar9__recorder_sn_vhold)) ;
assign post_value_holder_triggered__p191__ = (!(__IEND__))||((__auxvar10__recorder_sn_condmet)||(__auxvar10__recorder_sn_cond)) ;
assign post_value_holder_triggered__p192__ = (!(__IEND__))||((__auxvar11__recorder_sn_condmet)||(__auxvar11__recorder_sn_cond)) ;
assign post_value_holder_triggered__p193__ = (!(__IEND__))||((__auxvar12__recorder_sn_condmet)||(__auxvar12__recorder_sn_cond)) ;
assign post_value_holder_triggered__p194__ = (!(__IEND__))||((__auxvar13__recorder_sn_condmet)||(__auxvar13__recorder_sn_cond)) ;
assign post_value_holder_triggered__p195__ = (!(__IEND__))||((__auxvar14__recorder_sn_condmet)||(__auxvar14__recorder_sn_cond)) ;
assign post_value_holder_triggered__p196__ = (!(__IEND__))||((__auxvar15__recorder_sn_condmet)||(__auxvar15__recorder_sn_cond)) ;
assign post_value_holder_triggered__p197__ = (!(__IEND__))||((__auxvar16__recorder_sn_condmet)||(__auxvar16__recorder_sn_cond)) ;
assign post_value_holder_triggered__p198__ = (!(__IEND__))||((__auxvar17__recorder_sn_condmet)||(__auxvar17__recorder_sn_cond)) ;
assign post_value_holder_triggered__p199__ = (!(__IEND__))||((__auxvar18__recorder_sn_condmet)||(__auxvar18__recorder_sn_cond)) ;
assign post_value_holder_triggered__p200__ = (!(__IEND__))||((__auxvar19__recorder_sn_condmet)||(__auxvar19__recorder_sn_cond)) ;
assign post_value_holder_triggered__p201__ = (!(__IEND__))||((__auxvar1__recorder_sn_condmet)||(__auxvar1__recorder_sn_cond)) ;
assign post_value_holder_triggered__p202__ = (!(__IEND__))||((__auxvar20__recorder_sn_condmet)||(__auxvar20__recorder_sn_cond)) ;
assign post_value_holder_triggered__p203__ = (!(__IEND__))||((__auxvar21__recorder_sn_condmet)||(__auxvar21__recorder_sn_cond)) ;
assign post_value_holder_triggered__p204__ = (!(__IEND__))||((__auxvar22__recorder_sn_condmet)||(__auxvar22__recorder_sn_cond)) ;
assign post_value_holder_triggered__p205__ = (!(__IEND__))||((__auxvar23__recorder_sn_condmet)||(__auxvar23__recorder_sn_cond)) ;
assign post_value_holder_triggered__p206__ = (!(__IEND__))||((__auxvar24__recorder_sn_condmet)||(__auxvar24__recorder_sn_cond)) ;
assign post_value_holder_triggered__p207__ = (!(__IEND__))||((__auxvar25__recorder_sn_condmet)||(__auxvar25__recorder_sn_cond)) ;
assign post_value_holder_triggered__p208__ = (!(__IEND__))||((__auxvar26__recorder_sn_condmet)||(__auxvar26__recorder_sn_cond)) ;
assign post_value_holder_triggered__p209__ = (!(__IEND__))||((__auxvar27__recorder_sn_condmet)||(__auxvar27__recorder_sn_cond)) ;
assign post_value_holder_triggered__p210__ = (!(__IEND__))||((__auxvar28__recorder_sn_condmet)||(__auxvar28__recorder_sn_cond)) ;
assign post_value_holder_triggered__p211__ = (!(__IEND__))||((__auxvar29__recorder_sn_condmet)||(__auxvar29__recorder_sn_cond)) ;
assign post_value_holder_triggered__p212__ = (!(__IEND__))||((__auxvar2__recorder_sn_condmet)||(__auxvar2__recorder_sn_cond)) ;
assign post_value_holder_triggered__p213__ = (!(__IEND__))||((__auxvar30__recorder_sn_condmet)||(__auxvar30__recorder_sn_cond)) ;
assign post_value_holder_triggered__p214__ = (!(__IEND__))||((__auxvar31__recorder_sn_condmet)||(__auxvar31__recorder_sn_cond)) ;
assign post_value_holder_triggered__p215__ = (!(__IEND__))||((__auxvar32__recorder_sn_condmet)||(__auxvar32__recorder_sn_cond)) ;
assign post_value_holder_triggered__p216__ = (!(__IEND__))||((__auxvar33__recorder_sn_condmet)||(__auxvar33__recorder_sn_cond)) ;
assign post_value_holder_triggered__p217__ = (!(__IEND__))||((__auxvar34__recorder_sn_condmet)||(__auxvar34__recorder_sn_cond)) ;
assign post_value_holder_triggered__p218__ = (!(__IEND__))||((__auxvar35__recorder_sn_condmet)||(__auxvar35__recorder_sn_cond)) ;
assign post_value_holder_triggered__p219__ = (!(__IEND__))||((__auxvar36__recorder_sn_condmet)||(__auxvar36__recorder_sn_cond)) ;
assign post_value_holder_triggered__p220__ = (!(__IEND__))||((__auxvar37__recorder_sn_condmet)||(__auxvar37__recorder_sn_cond)) ;
assign post_value_holder_triggered__p221__ = (!(__IEND__))||((__auxvar38__recorder_sn_condmet)||(__auxvar38__recorder_sn_cond)) ;
assign post_value_holder_triggered__p222__ = (!(__IEND__))||((__auxvar3__recorder_sn_condmet)||(__auxvar3__recorder_sn_cond)) ;
assign post_value_holder_triggered__p223__ = (!(__IEND__))||((__auxvar4__recorder_sn_condmet)||(__auxvar4__recorder_sn_cond)) ;
assign post_value_holder_triggered__p224__ = (!(__IEND__))||((__auxvar5__recorder_sn_condmet)||(__auxvar5__recorder_sn_cond)) ;
assign post_value_holder_triggered__p225__ = (!(__IEND__))||((__auxvar6__recorder_sn_condmet)||(__auxvar6__recorder_sn_cond)) ;
assign post_value_holder_triggered__p226__ = (!(__IEND__))||((__auxvar7__recorder_sn_condmet)||(__auxvar7__recorder_sn_cond)) ;
assign post_value_holder_triggered__p227__ = (!(__IEND__))||((__auxvar8__recorder_sn_condmet)||(__auxvar8__recorder_sn_cond)) ;
assign post_value_holder_triggered__p228__ = (!(__IEND__))||((__auxvar9__recorder_sn_condmet)||(__auxvar9__recorder_sn_cond)) ;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem$dmem_req_op;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL__RTL__DOT__rg_trap_instr;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire[63:0] RTL__RTL__DOT__near_mem$dmem_req_store_value;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire[63:0] RTL__RTL__DOT__near_mem$dmem_word64;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    wire[31:0] RTL__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__RTL__DOT__s1_to_s2$D_IN;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    wire RTL__RTL__DOT__stage2_rg_full;
    wire RTL__RTL__DOT__csr_regfile__DOT__rg_state;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__RTL__DOT__stage1_rg_full;
    wire RTL__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    wire RTL__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL__RTL__DOT__rg_run_on_reset;
    wire RTL__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL__RTL__DOT__s2_to_s3$EN;
    wire[2:0] RTL__RTL__DOT__near_mem$dmem_req_f3;
    wire RTL__RTL__DOT__s1_to_s2$EN;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    wire RTL__RTL__DOT__s3_deq$EN;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire[3:0] RTL__RTL__DOT__rg_state;
    wire RTL__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__RTL__DOT__rg_retiring$EN;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__RTL__DOT__s2_to_s3$D_IN;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    wire RTL__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL__RTL__DOT__stage3_rg_full;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    wire[168:0] RTL__RTL__DOT__stage2_rg_stage2;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    wire RTL__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__RTL__DOT__csr_regfile__DOT__rg_nmi;
    wire[31:0] RTL__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL__RTL__DOT__near_mem$EN_dmem_req;
    wire RTL__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire[1:0] RTL__RTL__DOT__rg_cur_priv;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    wire RTL__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    wire[31:0] RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire[31:0] RTL__RTL__DOT__near_mem$dmem_req_addr;
    wire[31:0] RTL__RTL__DOT__near_mem$imem_instr;
    wire RTL__RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire[31:0] RTL__RTL__DOT__near_mem$imem_pc;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem$dmem_exc;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__RTL__DOT__s3_deq$D_IN;
    wire RTL__CLK;
    wire RTL__RST_N;
    wire RTL__hart0_server_reset_request_put;
    wire RTL__EN_hart0_server_reset_request_put;
    wire RTL__RDY_hart0_server_reset_request_put;
    wire RTL__EN_hart0_server_reset_response_get;
    wire RTL__hart0_server_reset_response_get;
    wire RTL__RDY_hart0_server_reset_response_get;
    wire RTL__imem_master_awvalid;
    wire[3:0] RTL__imem_master_awid;
    wire[63:0] RTL__imem_master_awaddr;
    wire[7:0] RTL__imem_master_awlen;
    wire[2:0] RTL__imem_master_awsize;
    wire[1:0] RTL__imem_master_awburst;
    wire RTL__imem_master_awlock;
    wire[3:0] RTL__imem_master_awcache;
    wire[2:0] RTL__imem_master_awprot;
    wire[3:0] RTL__imem_master_awqos;
    wire[3:0] RTL__imem_master_awregion;
    wire RTL__imem_master_awready;
    wire RTL__imem_master_wvalid;
    wire[63:0] RTL__imem_master_wdata;
    wire[7:0] RTL__imem_master_wstrb;
    wire RTL__imem_master_wlast;
    wire RTL__imem_master_wready;
    wire RTL__imem_master_bvalid;
    wire[3:0] RTL__imem_master_bid;
    wire[1:0] RTL__imem_master_bresp;
    wire RTL__imem_master_bready;
    wire RTL__imem_master_arvalid;
    wire[3:0] RTL__imem_master_arid;
    wire[63:0] RTL__imem_master_araddr;
    wire[7:0] RTL__imem_master_arlen;
    wire[2:0] RTL__imem_master_arsize;
    wire[1:0] RTL__imem_master_arburst;
    wire RTL__imem_master_arlock;
    wire[3:0] RTL__imem_master_arcache;
    wire[2:0] RTL__imem_master_arprot;
    wire[3:0] RTL__imem_master_arqos;
    wire[3:0] RTL__imem_master_arregion;
    wire RTL__imem_master_arready;
    wire RTL__imem_master_rvalid;
    wire[3:0] RTL__imem_master_rid;
    wire[63:0] RTL__imem_master_rdata;
    wire[1:0] RTL__imem_master_rresp;
    wire RTL__imem_master_rlast;
    wire RTL__imem_master_rready;
    wire RTL__dmem_master_awvalid;
    wire[3:0] RTL__dmem_master_awid;
    wire[63:0] RTL__dmem_master_awaddr;
    wire[7:0] RTL__dmem_master_awlen;
    wire[2:0] RTL__dmem_master_awsize;
    wire[1:0] RTL__dmem_master_awburst;
    wire RTL__dmem_master_awlock;
    wire[3:0] RTL__dmem_master_awcache;
    wire[2:0] RTL__dmem_master_awprot;
    wire[3:0] RTL__dmem_master_awqos;
    wire[3:0] RTL__dmem_master_awregion;
    wire RTL__dmem_master_awready;
    wire RTL__dmem_master_wvalid;
    wire[63:0] RTL__dmem_master_wdata;
    wire[7:0] RTL__dmem_master_wstrb;
    wire RTL__dmem_master_wlast;
    wire RTL__dmem_master_wready;
    wire RTL__dmem_master_bvalid;
    wire[3:0] RTL__dmem_master_bid;
    wire[1:0] RTL__dmem_master_bresp;
    wire RTL__dmem_master_bready;
    wire RTL__dmem_master_arvalid;
    wire[3:0] RTL__dmem_master_arid;
    wire[63:0] RTL__dmem_master_araddr;
    wire[7:0] RTL__dmem_master_arlen;
    wire[2:0] RTL__dmem_master_arsize;
    wire[1:0] RTL__dmem_master_arburst;
    wire RTL__dmem_master_arlock;
    wire[3:0] RTL__dmem_master_arcache;
    wire[2:0] RTL__dmem_master_arprot;
    wire[3:0] RTL__dmem_master_arqos;
    wire[3:0] RTL__dmem_master_arregion;
    wire RTL__dmem_master_arready;
    wire RTL__dmem_master_rvalid;
    wire[3:0] RTL__dmem_master_rid;
    wire[63:0] RTL__dmem_master_rdata;
    wire[1:0] RTL__dmem_master_rresp;
    wire RTL__dmem_master_rlast;
    wire RTL__dmem_master_rready;
    wire RTL__m_external_interrupt_req_set_not_clear;
    wire RTL__s_external_interrupt_req_set_not_clear;
    wire RTL__software_interrupt_req_set_not_clear;
    wire RTL__timer_interrupt_req_set_not_clear;
    wire RTL__nmi_req_set_not_clear;
    wire[3:0] RTL__set_verbosity_verbosity;
    wire[63:0] RTL__set_verbosity_logdelay;
    wire RTL__EN_set_verbosity;
    wire RTL__RDY_set_verbosity;

    wire[63:0] RTL__dmem_master_araddr , RTL__dmem_master_awaddr , RTL__dmem_master_wdata , RTL__imem_master_araddr , RTL__imem_master_awaddr , RTL__imem_master_wdata ; 
    wire[7:0] RTL__dmem_master_arlen , RTL__dmem_master_awlen , RTL__dmem_master_wstrb , RTL__imem_master_arlen , RTL__imem_master_awlen , RTL__imem_master_wstrb ; 
    wire[3:0] RTL__dmem_master_arcache , RTL__dmem_master_arid , RTL__dmem_master_arqos , RTL__dmem_master_arregion , RTL__dmem_master_awcache , RTL__dmem_master_awid , RTL__dmem_master_awqos , RTL__dmem_master_awregion , RTL__imem_master_arcache , RTL__imem_master_arid , RTL__imem_master_arqos , RTL__imem_master_arregion , RTL__imem_master_awcache , RTL__imem_master_awid , RTL__imem_master_awqos , RTL__imem_master_awregion ; 
    wire[2:0] RTL__dmem_master_arprot , RTL__dmem_master_arsize , RTL__dmem_master_awprot , RTL__dmem_master_awsize , RTL__imem_master_arprot , RTL__imem_master_arsize , RTL__imem_master_awprot , RTL__imem_master_awsize ; 
    wire[1:0] RTL__dmem_master_arburst , RTL__dmem_master_awburst , RTL__imem_master_arburst , RTL__imem_master_awburst ; 
    wire RTL__RDY_hart0_server_reset_request_put , RTL__RDY_hart0_server_reset_response_get , RTL__RDY_set_verbosity , RTL__dmem_master_arlock , RTL__dmem_master_arvalid , RTL__dmem_master_awlock , RTL__dmem_master_awvalid , RTL__dmem_master_bready , RTL__dmem_master_rready , RTL__dmem_master_wlast , RTL__dmem_master_wvalid , RTL__hart0_server_reset_response_get , RTL__imem_master_arlock , RTL__imem_master_arvalid , RTL__imem_master_awlock , RTL__imem_master_awvalid , RTL__imem_master_bready , RTL__imem_master_rready , RTL__imem_master_wlast , RTL__imem_master_wvalid ; reg[63:0] RTL__cfg_logdelay ; 
    wire[63:0] RTL__cfg_logdelay$D_IN ; 
    wire RTL__cfg_logdelay$EN ; reg[3:0] RTL__cfg_verbosity ; 
    wire[3:0] RTL__cfg_verbosity$D_IN ; 
    wire RTL__cfg_verbosity$EN ; reg[31:0] RTL__rg_csr_pc ; 
    wire[31:0] RTL__rg_csr_pc$D_IN ; 
    wire RTL__rg_csr_pc$EN ; reg[31:0] RTL__rg_csr_val1 ; 
    wire[31:0] RTL__rg_csr_val1$D_IN ; 
    wire RTL__rg_csr_val1$EN ; reg[1:0] RTL__rg_cur_priv ; reg[1:0] RTL__rg_cur_priv$D_IN ; 
    wire RTL__rg_cur_priv$EN ; 
    reg RTL__rg_mstatus_MXR ; 
    wire RTL__rg_mstatus_MXR$D_IN , RTL__rg_mstatus_MXR$EN ; reg[31:0] RTL__rg_next_pc ; reg[31:0] RTL__rg_next_pc$D_IN ; 
    wire RTL__rg_next_pc$EN ; 
    reg RTL__rg_retiring ; 
    wire RTL__rg_retiring$D_IN , RTL__rg_retiring$EN ; 
    reg RTL__rg_run_on_reset ; 
    wire RTL__rg_run_on_reset$D_IN , RTL__rg_run_on_reset$EN ; 
    reg RTL__rg_sstatus_SUM ; 
    wire RTL__rg_sstatus_SUM$D_IN , RTL__rg_sstatus_SUM$EN ; reg[63:0] RTL__rg_start_CPI_cycles ; 
    wire[63:0] RTL__rg_start_CPI_cycles$D_IN ; 
    wire RTL__rg_start_CPI_cycles$EN ; reg[63:0] RTL__rg_start_CPI_instrs ; 
    wire[63:0] RTL__rg_start_CPI_instrs$D_IN ; 
    wire RTL__rg_start_CPI_instrs$EN ; reg[3:0] RTL__rg_state ; reg[3:0] RTL__rg_state$D_IN ; 
    wire RTL__rg_state$EN ; reg[67:0] RTL__rg_trap_info ; reg[67:0] RTL__rg_trap_info$D_IN ; 
    wire RTL__rg_trap_info$EN ; reg[31:0] RTL__rg_trap_instr ; 
    wire[31:0] RTL__rg_trap_instr$D_IN ; 
    wire RTL__rg_trap_instr$EN ; 
    reg RTL__rg_trap_interrupt ; 
    wire RTL__rg_trap_interrupt$D_IN , RTL__rg_trap_interrupt$EN ; 
    reg RTL__s1_to_s2 ; 
    wire RTL__s1_to_s2$D_IN , RTL__s1_to_s2$EN ; 
    reg RTL__s2_to_s3 ; 
    wire RTL__s2_to_s3$D_IN , RTL__s2_to_s3$EN ; 
    reg RTL__s3_deq ; 
    wire RTL__s3_deq$D_IN , RTL__s3_deq$EN ; 
    reg RTL__stage1_rg_full ; 
    reg RTL__stage1_rg_full$D_IN ; 
    wire RTL__stage1_rg_full$EN ; 
    reg RTL__stage2_rg_full ; 
    reg RTL__stage2_rg_full$D_IN ; 
    wire RTL__stage2_rg_full$EN ; 
    reg RTL__stage2_rg_resetting ; 
    wire RTL__stage2_rg_resetting$D_IN , RTL__stage2_rg_resetting$EN ; reg[168:0] RTL__stage2_rg_stage2 ; 
    wire[168:0] RTL__stage2_rg_stage2$D_IN ; 
    wire RTL__stage2_rg_stage2$EN ; 
    reg RTL__stage3_rg_full ; 
    reg RTL__stage3_rg_full$D_IN ; 
    wire RTL__stage3_rg_full$EN ; reg[103:0] RTL__stage3_rg_stage3 ; 
    wire[103:0] RTL__stage3_rg_stage3$D_IN ; 
    wire RTL__stage3_rg_stage3$EN ; reg[1:0] RTL__csr_regfile$csr_ret_actions_from_priv ; 
    wire[97:0] RTL__csr_regfile$csr_trap_actions ; 
    wire[65:0] RTL__csr_regfile$csr_ret_actions ; 
    wire[63:0] RTL__csr_regfile$read_csr_mcycle , RTL__csr_regfile$read_csr_minstret ; 
    wire[32:0] RTL__csr_regfile$read_csr ; 
    wire[31:0] RTL__csr_regfile$csr_trap_actions_pc , RTL__csr_regfile$csr_trap_actions_xtval , RTL__csr_regfile$mav_csr_write_word , RTL__csr_regfile$read_mstatus , RTL__csr_regfile$read_satp ; 
    wire[27:0] RTL__csr_regfile$read_misa ; 
    wire[11:0] RTL__csr_regfile$access_permitted_1_csr_addr , RTL__csr_regfile$access_permitted_2_csr_addr , RTL__csr_regfile$csr_counter_read_fault_csr_addr , RTL__csr_regfile$mav_csr_write_csr_addr , RTL__csr_regfile$mav_read_csr_csr_addr , RTL__csr_regfile$read_csr_csr_addr , RTL__csr_regfile$read_csr_port2_csr_addr ; 
    wire[4:0] RTL__csr_regfile$interrupt_pending ; 
    wire[3:0] RTL__csr_regfile$csr_trap_actions_exc_code ; 
    wire[1:0] RTL__csr_regfile$access_permitted_1_priv , RTL__csr_regfile$access_permitted_2_priv , RTL__csr_regfile$csr_counter_read_fault_priv , RTL__csr_regfile$csr_trap_actions_from_priv , RTL__csr_regfile$interrupt_pending_cur_priv ; 
    wire RTL__csr_regfile$EN_csr_minstret_incr , RTL__csr_regfile$EN_csr_ret_actions , RTL__csr_regfile$EN_csr_trap_actions , RTL__csr_regfile$EN_debug , RTL__csr_regfile$EN_mav_csr_write , RTL__csr_regfile$EN_mav_read_csr , RTL__csr_regfile$EN_server_reset_request_put , RTL__csr_regfile$EN_server_reset_response_get , RTL__csr_regfile$RDY_server_reset_request_put , RTL__csr_regfile$RDY_server_reset_response_get , RTL__csr_regfile$access_permitted_1 , RTL__csr_regfile$access_permitted_1_read_not_write , RTL__csr_regfile$access_permitted_2 , RTL__csr_regfile$access_permitted_2_read_not_write , RTL__csr_regfile$csr_trap_actions_interrupt , RTL__csr_regfile$csr_trap_actions_nmi , RTL__csr_regfile$m_external_interrupt_req_set_not_clear , RTL__csr_regfile$nmi_pending , RTL__csr_regfile$nmi_req_set_not_clear , RTL__csr_regfile$s_external_interrupt_req_set_not_clear , RTL__csr_regfile$software_interrupt_req_set_not_clear , RTL__csr_regfile$timer_interrupt_req_set_not_clear , RTL__csr_regfile$wfi_resume ; 
    wire RTL__f_reset_reqs$CLR , RTL__f_reset_reqs$DEQ , RTL__f_reset_reqs$D_IN , RTL__f_reset_reqs$D_OUT , RTL__f_reset_reqs$EMPTY_N , RTL__f_reset_reqs$ENQ , RTL__f_reset_reqs$FULL_N ; 
    wire RTL__f_reset_rsps$CLR , RTL__f_reset_rsps$DEQ , RTL__f_reset_rsps$D_IN , RTL__f_reset_rsps$D_OUT , RTL__f_reset_rsps$EMPTY_N , RTL__f_reset_rsps$ENQ , RTL__f_reset_rsps$FULL_N ; 
    wire[31:0] RTL__gpr_regfile$read_rs1 , RTL__gpr_regfile$read_rs2 , RTL__gpr_regfile$write_rd_rd_val ; 
    wire[4:0] RTL__gpr_regfile$read_rs1_port2_rs1 , RTL__gpr_regfile$read_rs1_rs1 , RTL__gpr_regfile$read_rs2_rs2 , RTL__gpr_regfile$write_rd_rd ; 
    wire RTL__gpr_regfile$EN_server_reset_request_put , RTL__gpr_regfile$EN_server_reset_response_get , RTL__gpr_regfile$EN_write_rd , RTL__gpr_regfile$RDY_server_reset_request_put , RTL__gpr_regfile$RDY_server_reset_response_get ; reg[31:0] RTL__near_mem$imem_req_addr ; 
    wire[63:0] RTL__near_mem$dmem_master_araddr , RTL__near_mem$dmem_master_awaddr , RTL__near_mem$dmem_master_rdata , RTL__near_mem$dmem_master_wdata , RTL__near_mem$dmem_req_store_value , RTL__near_mem$dmem_word64 , RTL__near_mem$imem_master_araddr , RTL__near_mem$imem_master_awaddr , RTL__near_mem$imem_master_rdata , RTL__near_mem$imem_master_wdata ; 
    wire[31:0] RTL__near_mem$dmem_req_addr , RTL__near_mem$dmem_req_satp , RTL__near_mem$imem_instr , RTL__near_mem$imem_pc , RTL__near_mem$imem_req_satp , RTL__near_mem$imem_tval ; 
    wire[7:0] RTL__near_mem$dmem_master_arlen , RTL__near_mem$dmem_master_awlen , RTL__near_mem$dmem_master_wstrb , RTL__near_mem$imem_master_arlen , RTL__near_mem$imem_master_awlen , RTL__near_mem$imem_master_wstrb , RTL__near_mem$server_fence_request_put ; 
    wire[3:0] RTL__near_mem$dmem_exc_code , RTL__near_mem$dmem_master_arcache , RTL__near_mem$dmem_master_arid , RTL__near_mem$dmem_master_arqos , RTL__near_mem$dmem_master_arregion , RTL__near_mem$dmem_master_awcache , RTL__near_mem$dmem_master_awid , RTL__near_mem$dmem_master_awqos , RTL__near_mem$dmem_master_awregion , RTL__near_mem$dmem_master_bid , RTL__near_mem$dmem_master_rid , RTL__near_mem$imem_exc_code , RTL__near_mem$imem_master_arcache , RTL__near_mem$imem_master_arid , RTL__near_mem$imem_master_arqos , RTL__near_mem$imem_master_arregion , RTL__near_mem$imem_master_awcache , RTL__near_mem$imem_master_awid , RTL__near_mem$imem_master_awqos , RTL__near_mem$imem_master_awregion , RTL__near_mem$imem_master_bid , RTL__near_mem$imem_master_rid ; 
    wire[2:0] RTL__near_mem$dmem_master_arprot , RTL__near_mem$dmem_master_arsize , RTL__near_mem$dmem_master_awprot , RTL__near_mem$dmem_master_awsize , RTL__near_mem$dmem_req_f3 , RTL__near_mem$imem_master_arprot , RTL__near_mem$imem_master_arsize , RTL__near_mem$imem_master_awprot , RTL__near_mem$imem_master_awsize , RTL__near_mem$imem_req_f3 ; 
    wire[1:0] RTL__near_mem$dmem_master_arburst , RTL__near_mem$dmem_master_awburst , RTL__near_mem$dmem_master_bresp , RTL__near_mem$dmem_master_rresp , RTL__near_mem$dmem_req_priv , RTL__near_mem$imem_master_arburst , RTL__near_mem$imem_master_awburst , RTL__near_mem$imem_master_bresp , RTL__near_mem$imem_master_rresp , RTL__near_mem$imem_req_priv ; 
    wire RTL__near_mem$EN_dmem_req , RTL__near_mem$EN_imem_req , RTL__near_mem$EN_server_fence_i_request_put , RTL__near_mem$EN_server_fence_i_response_get , RTL__near_mem$EN_server_fence_request_put , RTL__near_mem$EN_server_fence_response_get , RTL__near_mem$EN_server_reset_request_put , RTL__near_mem$EN_server_reset_response_get , RTL__near_mem$EN_sfence_vma , RTL__near_mem$RDY_server_fence_i_request_put , RTL__near_mem$RDY_server_fence_i_response_get , RTL__near_mem$RDY_server_fence_request_put , RTL__near_mem$RDY_server_fence_response_get , RTL__near_mem$RDY_server_reset_request_put , RTL__near_mem$RDY_server_reset_response_get , RTL__near_mem$dmem_exc , RTL__near_mem$dmem_master_arlock , RTL__near_mem$dmem_master_arready , RTL__near_mem$dmem_master_arvalid , RTL__near_mem$dmem_master_awlock , RTL__near_mem$dmem_master_awready , RTL__near_mem$dmem_master_awvalid , RTL__near_mem$dmem_master_bready , RTL__near_mem$dmem_master_bvalid , RTL__near_mem$dmem_master_rlast , RTL__near_mem$dmem_master_rready , RTL__near_mem$dmem_master_rvalid , RTL__near_mem$dmem_master_wlast , RTL__near_mem$dmem_master_wready , RTL__near_mem$dmem_master_wvalid , RTL__near_mem$dmem_req_mstatus_MXR , RTL__near_mem$dmem_req_op , RTL__near_mem$dmem_req_sstatus_SUM , RTL__near_mem$dmem_valid , RTL__near_mem$imem_exc , RTL__near_mem$imem_is_i32_not_i16 , RTL__near_mem$imem_master_arlock , RTL__near_mem$imem_master_arready , RTL__near_mem$imem_master_arvalid , RTL__near_mem$imem_master_awlock , RTL__near_mem$imem_master_awready , RTL__near_mem$imem_master_awvalid , RTL__near_mem$imem_master_bready , RTL__near_mem$imem_master_bvalid , RTL__near_mem$imem_master_rlast , RTL__near_mem$imem_master_rready , RTL__near_mem$imem_master_rvalid , RTL__near_mem$imem_master_wlast , RTL__near_mem$imem_master_wready , RTL__near_mem$imem_master_wvalid , RTL__near_mem$imem_req_mstatus_MXR , RTL__near_mem$imem_req_sstatus_SUM , RTL__near_mem$imem_valid ; 
    wire[63:0] RTL__soc_map$m_is_IO_addr_addr , RTL__soc_map$m_is_mem_addr_addr , RTL__soc_map$m_is_near_mem_IO_addr_addr , RTL__soc_map$m_pc_reset_value ; 
    wire RTL__stage1_f_reset_reqs$CLR , RTL__stage1_f_reset_reqs$DEQ , RTL__stage1_f_reset_reqs$EMPTY_N , RTL__stage1_f_reset_reqs$ENQ , RTL__stage1_f_reset_reqs$FULL_N ; 
    wire RTL__stage1_f_reset_rsps$CLR , RTL__stage1_f_reset_rsps$DEQ , RTL__stage1_f_reset_rsps$EMPTY_N , RTL__stage1_f_reset_rsps$ENQ , RTL__stage1_f_reset_rsps$FULL_N ; 
    wire RTL__stage2_f_reset_reqs$CLR , RTL__stage2_f_reset_reqs$DEQ , RTL__stage2_f_reset_reqs$EMPTY_N , RTL__stage2_f_reset_reqs$ENQ , RTL__stage2_f_reset_reqs$FULL_N ; 
    wire RTL__stage2_f_reset_rsps$CLR , RTL__stage2_f_reset_rsps$DEQ , RTL__stage2_f_reset_rsps$EMPTY_N , RTL__stage2_f_reset_rsps$ENQ , RTL__stage2_f_reset_rsps$FULL_N ; 
    wire RTL__stage3_f_reset_reqs$CLR , RTL__stage3_f_reset_reqs$DEQ , RTL__stage3_f_reset_reqs$EMPTY_N , RTL__stage3_f_reset_reqs$ENQ , RTL__stage3_f_reset_reqs$FULL_N ; 
    wire RTL__stage3_f_reset_rsps$CLR , RTL__stage3_f_reset_rsps$DEQ , RTL__stage3_f_reset_rsps$EMPTY_N , RTL__stage3_f_reset_rsps$ENQ , RTL__stage3_f_reset_rsps$FULL_N ; 
    wire RTL__CAN_FIRE_RL_rl_WFI_resume , RTL__CAN_FIRE_RL_rl_finish_FENCE , RTL__CAN_FIRE_RL_rl_finish_FENCE_I , RTL__CAN_FIRE_RL_rl_finish_SFENCE_VMA , RTL__CAN_FIRE_RL_rl_pipe , RTL__CAN_FIRE_RL_rl_reset_complete , RTL__CAN_FIRE_RL_rl_reset_from_WFI , RTL__CAN_FIRE_RL_rl_reset_start , RTL__CAN_FIRE_RL_rl_show_pipe , RTL__CAN_FIRE_RL_rl_stage1_CSRR_S_or_C , RTL__CAN_FIRE_RL_rl_stage1_CSRR_S_or_C_2 , RTL__CAN_FIRE_RL_rl_stage1_CSRR_W , RTL__CAN_FIRE_RL_rl_stage1_CSRR_W_2 , RTL__CAN_FIRE_RL_rl_stage1_FENCE , RTL__CAN_FIRE_RL_rl_stage1_FENCE_I , RTL__CAN_FIRE_RL_rl_stage1_SFENCE_VMA , RTL__CAN_FIRE_RL_rl_stage1_WFI , RTL__CAN_FIRE_RL_rl_stage1_interrupt , RTL__CAN_FIRE_RL_rl_stage1_restart_after_csrrx , RTL__CAN_FIRE_RL_rl_stage1_trap , RTL__CAN_FIRE_RL_rl_stage1_xRET , RTL__CAN_FIRE_RL_rl_stage2_nonpipe , RTL__CAN_FIRE_RL_rl_trap , RTL__CAN_FIRE_RL_rl_trap_fetch , RTL__CAN_FIRE_RL_stage1_rl_reset , RTL__CAN_FIRE_RL_stage2_rl_reset_begin , RTL__CAN_FIRE_RL_stage2_rl_reset_end , RTL__CAN_FIRE_RL_stage3_rl_reset , RTL__CAN_FIRE_dmem_master_m_arready , RTL__CAN_FIRE_dmem_master_m_awready , RTL__CAN_FIRE_dmem_master_m_bvalid , RTL__CAN_FIRE_dmem_master_m_rvalid , RTL__CAN_FIRE_dmem_master_m_wready , RTL__CAN_FIRE_hart0_server_reset_request_put , RTL__CAN_FIRE_hart0_server_reset_response_get , RTL__CAN_FIRE_imem_master_m_arready , RTL__CAN_FIRE_imem_master_m_awready , RTL__CAN_FIRE_imem_master_m_bvalid , RTL__CAN_FIRE_imem_master_m_rvalid , RTL__CAN_FIRE_imem_master_m_wready , RTL__CAN_FIRE_m_external_interrupt_req , RTL__CAN_FIRE_nmi_req , RTL__CAN_FIRE_s_external_interrupt_req , RTL__CAN_FIRE_set_verbosity , RTL__CAN_FIRE_software_interrupt_req , RTL__CAN_FIRE_timer_interrupt_req , RTL__WILL_FIRE_RL_rl_WFI_resume , RTL__WILL_FIRE_RL_rl_finish_FENCE , RTL__WILL_FIRE_RL_rl_finish_FENCE_I , RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA , RTL__WILL_FIRE_RL_rl_pipe , RTL__WILL_FIRE_RL_rl_reset_complete , RTL__WILL_FIRE_RL_rl_reset_from_WFI , RTL__WILL_FIRE_RL_rl_reset_start , RTL__WILL_FIRE_RL_rl_show_pipe , RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C , RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 , RTL__WILL_FIRE_RL_rl_stage1_CSRR_W , RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 , RTL__WILL_FIRE_RL_rl_stage1_FENCE , RTL__WILL_FIRE_RL_rl_stage1_FENCE_I , RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA , RTL__WILL_FIRE_RL_rl_stage1_WFI , RTL__WILL_FIRE_RL_rl_stage1_interrupt , RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx , RTL__WILL_FIRE_RL_rl_stage1_trap , RTL__WILL_FIRE_RL_rl_stage1_xRET , RTL__WILL_FIRE_RL_rl_stage2_nonpipe , RTL__WILL_FIRE_RL_rl_trap , RTL__WILL_FIRE_RL_rl_trap_fetch , RTL__WILL_FIRE_RL_stage1_rl_reset , RTL__WILL_FIRE_RL_stage2_rl_reset_begin , RTL__WILL_FIRE_RL_stage2_rl_reset_end , RTL__WILL_FIRE_RL_stage3_rl_reset , RTL__WILL_FIRE_dmem_master_m_arready , RTL__WILL_FIRE_dmem_master_m_awready , RTL__WILL_FIRE_dmem_master_m_bvalid , RTL__WILL_FIRE_dmem_master_m_rvalid , RTL__WILL_FIRE_dmem_master_m_wready , RTL__WILL_FIRE_hart0_server_reset_request_put , RTL__WILL_FIRE_hart0_server_reset_response_get , RTL__WILL_FIRE_imem_master_m_arready , RTL__WILL_FIRE_imem_master_m_awready , RTL__WILL_FIRE_imem_master_m_bvalid , RTL__WILL_FIRE_imem_master_m_rvalid , RTL__WILL_FIRE_imem_master_m_wready , RTL__WILL_FIRE_m_external_interrupt_req , RTL__WILL_FIRE_nmi_req , RTL__WILL_FIRE_s_external_interrupt_req , RTL__WILL_FIRE_set_verbosity , RTL__WILL_FIRE_software_interrupt_req , RTL__WILL_FIRE_timer_interrupt_req ; reg[31:0] RTL__MUX_csr_regfile$mav_csr_write_2__VAL_2 ; 
    wire[67:0] RTL__MUX_rg_trap_info$write_1__VAL_1 , RTL__MUX_rg_trap_info$write_1__VAL_2 , RTL__MUX_rg_trap_info$write_1__VAL_3 , RTL__MUX_rg_trap_info$write_1__VAL_4 ; 
    wire[3:0] RTL__MUX_rg_state$write_1__VAL_1 , RTL__MUX_rg_state$write_1__VAL_2 , RTL__MUX_rg_state$write_1__VAL_3 ; 
    wire RTL__MUX_csr_regfile$mav_csr_write_1__SEL_1 , RTL__MUX_gpr_regfile$write_rd_1__SEL_3 , RTL__MUX_near_mem$imem_req_1__SEL_1 , RTL__MUX_near_mem$imem_req_1__SEL_2 , RTL__MUX_near_mem$imem_req_1__SEL_5 , RTL__MUX_rg_next_pc$write_1__SEL_1 , RTL__MUX_rg_retiring$write_1__SEL_1 , RTL__MUX_rg_state$write_1__SEL_1 , RTL__MUX_rg_state$write_1__SEL_10 , RTL__MUX_rg_state$write_1__SEL_4 , RTL__MUX_rg_state$write_1__SEL_6 , RTL__MUX_rg_state$write_1__SEL_7 , RTL__MUX_rg_state$write_1__SEL_8 , RTL__MUX_rg_state$write_1__SEL_9 , RTL__MUX_rg_trap_info$write_1__SEL_1 , RTL__MUX_rg_trap_instr$write_1__SEL_1 , RTL__MUX_rg_trap_interrupt$write_1__SEL_1 , RTL__MUX_s1_to_s2$write_1__VAL_1 , RTL__MUX_stage1_rg_full$write_1__VAL_10 , RTL__MUX_stage2_rg_full$write_1__VAL_3 ; reg[31:0] RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570 , RTL___theResult_____1_fst__h6569 , RTL__rs1_val__h11920 , RTL__x_out_data_to_stage2_addr__h5223 , RTL__x_out_data_to_stage2_val1__h5224 , RTL__x_out_data_to_stage3_rd_val__h4668 ; reg[4:0] RTL__x_out_data_to_stage3_rd__h4667 ; reg[3:0] RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10 , RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12 , RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11 , RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13 , RTL__CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4 , RTL__CASE_rg_cur_priv_0b0_8_0b1_9_11__q3 , RTL__IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413 , RTL__alu_outputs_exc_code__h5862 ; reg[1:0] RTL__CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5 , RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ; 
    reg RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8 , RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9 , RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 , RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ; 
    wire[127:0] RTL__csr_regfile_read_csr_mcycle__8_MINUS_rg_start__ETC___d818 ; 
    wire[63:0] RTL___theResult____h10743 , RTL__cpi__h10745 , RTL__cpifrac__h10746 , RTL__delta_CPI_cycles__h10741 , RTL__delta_CPI_instrs___1__h10778 , RTL__delta_CPI_instrs__h10742 , RTL__x__h10744 ; 
    wire[35:0] RTL__IF_near_mem_imem_exc__78_THEN_near_mem_imem_ex_ETC___d799 ; 
    wire[31:0] RTL__IF_IF_near_mem_imem_instr__59_BITS_6_TO_0_79_E_ETC___d655 , RTL__IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571 , RTL__SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 , RTL___theResult_____1_fst__h6562 , RTL___theResult_____1_fst__h6597 , RTL___theResult___snd__h7382 , RTL__alu_outputs___1_addr__h5365 , RTL__alu_outputs___1_addr__h5385 , RTL__alu_outputs___1_addr__h5410 , RTL__alu_outputs___1_addr__h5583 , RTL__alu_outputs___1_val1__h5386 , RTL__alu_outputs___1_val1__h5480 , RTL__alu_outputs___1_val1__h5516 , RTL__alu_outputs___1_val1__h5847 , RTL__alu_outputs___1_val2__h5367 , RTL__data_to_stage2_addr__h5215 , RTL__eaddr__h5553 , RTL__fall_through_pc__h5175 , RTL__output_stage2___1_bypass_rd_val__h4960 , RTL__rd_val___1__h6550 , RTL__rd_val___1__h6558 , RTL__rd_val___1__h6565 , RTL__rd_val___1__h6572 , RTL__rd_val___1__h6579 , RTL__rd_val___1__h6586 , RTL__rd_val__h5072 , RTL__rd_val__h5132 , RTL__rd_val__h5523 , RTL__rd_val__h5537 , RTL__rd_val__h7278 , RTL__rd_val__h7330 , RTL__rd_val__h7352 , RTL__rs1_val__h11213 , RTL__rs1_val_bypassed__h3337 , RTL__rs2_val__h5339 , RTL__trap_info_tval__h6925 , RTL__val__h5074 , RTL__val__h5134 , RTL__value__h6967 , RTL__x_out_bypass_rd_val__h4969 , RTL__x_out_data_to_stage2_val2__h5225 , RTL__x_out_next_pc__h5189 , RTL__y__h12191 ; 
    wire[20:0] RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 ; 
    wire[12:0] RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 ; 
    wire[11:0] RTL__near_memimem_instr_BITS_31_TO_20__q7 , RTL__near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 ; 
    wire[4:0] RTL__shamt__h5467 , RTL__x_out_data_to_stage2_rd__h5222 ; 
    wire[3:0] RTL__IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362 , RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 , RTL__IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394 , RTL__alu_outputs___1_exc_code__h5362 , RTL__alu_outputs___1_exc_code__h5843 , RTL__cur_verbosity__h1827 , RTL__x_exc_code__h15410 , RTL__x_out_trap_info_exc_code__h6928 ; 
    wire[1:0] RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 , RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 , RTL__IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137 , RTL__IF_stage2_rg_stage2_4_BITS_102_TO_101_5_EQ_0_6_ETC___d85 ; 
    wire RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285 , RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 , RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 , RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d649 , RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d910 , RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 , RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 , RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 , RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d730 , RTL__NOT_IF_stage2_rg_full_3_THEN_IF_stage2_rg_stag_ETC___d109 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d769 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d776 , RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d790 , RTL__NOT_near_mem_imem_exc__78_13_AND_IF_near_mem_i_ETC___d481 , RTL__NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252 , RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 , RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 , RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 , RTL___0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 , RTL__csr_regfile_interrupt_pending_rg_cur_priv_9_07_ETC___d779 , RTL__gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 , RTL__gpr_regfile_RDY_server_reset_response_get__76__ETC___d688 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d578 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d581 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d584 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d587 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d590 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d593 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d596 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d599 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d602 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d605 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d608 , RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d611 , RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328 , RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616 , RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 , RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 , RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 , RTL__rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_EQ_0_ETC___d392 , RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 , RTL__rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 ; 
  assign  RTL__RDY_hart0_server_reset_request_put = RTL__f_reset_reqs$FULL_N ; 
  assign  RTL__CAN_FIRE_hart0_server_reset_request_put = RTL__f_reset_reqs$FULL_N ; 
  assign  RTL__WILL_FIRE_hart0_server_reset_request_put = RTL__EN_hart0_server_reset_request_put ; 
  assign  RTL__hart0_server_reset_response_get = RTL__f_reset_rsps$D_OUT ; 
  assign  RTL__RDY_hart0_server_reset_response_get = RTL__f_reset_rsps$EMPTY_N ; 
  assign  RTL__CAN_FIRE_hart0_server_reset_response_get = RTL__f_reset_rsps$EMPTY_N ; 
  assign  RTL__WILL_FIRE_hart0_server_reset_response_get = RTL__EN_hart0_server_reset_response_get ; 
  assign  RTL__imem_master_awvalid = RTL__near_mem$imem_master_awvalid ; 
  assign  RTL__imem_master_awid = RTL__near_mem$imem_master_awid ; 
  assign  RTL__imem_master_awaddr = RTL__near_mem$imem_master_awaddr ; 
  assign  RTL__imem_master_awlen = RTL__near_mem$imem_master_awlen ; 
  assign  RTL__imem_master_awsize = RTL__near_mem$imem_master_awsize ; 
  assign  RTL__imem_master_awburst = RTL__near_mem$imem_master_awburst ; 
  assign  RTL__imem_master_awlock = RTL__near_mem$imem_master_awlock ; 
  assign  RTL__imem_master_awcache = RTL__near_mem$imem_master_awcache ; 
  assign  RTL__imem_master_awprot = RTL__near_mem$imem_master_awprot ; 
  assign  RTL__imem_master_awqos = RTL__near_mem$imem_master_awqos ; 
  assign  RTL__imem_master_awregion = RTL__near_mem$imem_master_awregion ; 
  assign  RTL__CAN_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL__WILL_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL__imem_master_wvalid = RTL__near_mem$imem_master_wvalid ; 
  assign  RTL__imem_master_wdata = RTL__near_mem$imem_master_wdata ; 
  assign  RTL__imem_master_wstrb = RTL__near_mem$imem_master_wstrb ; 
  assign  RTL__imem_master_wlast = RTL__near_mem$imem_master_wlast ; 
  assign  RTL__CAN_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL__WILL_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL__CAN_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL__WILL_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL__imem_master_bready = RTL__near_mem$imem_master_bready ; 
  assign  RTL__imem_master_arvalid = RTL__near_mem$imem_master_arvalid ; 
  assign  RTL__imem_master_arid = RTL__near_mem$imem_master_arid ; 
  assign  RTL__imem_master_araddr = RTL__near_mem$imem_master_araddr ; 
  assign  RTL__imem_master_arlen = RTL__near_mem$imem_master_arlen ; 
  assign  RTL__imem_master_arsize = RTL__near_mem$imem_master_arsize ; 
  assign  RTL__imem_master_arburst = RTL__near_mem$imem_master_arburst ; 
  assign  RTL__imem_master_arlock = RTL__near_mem$imem_master_arlock ; 
  assign  RTL__imem_master_arcache = RTL__near_mem$imem_master_arcache ; 
  assign  RTL__imem_master_arprot = RTL__near_mem$imem_master_arprot ; 
  assign  RTL__imem_master_arqos = RTL__near_mem$imem_master_arqos ; 
  assign  RTL__imem_master_arregion = RTL__near_mem$imem_master_arregion ; 
  assign  RTL__CAN_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL__WILL_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL__CAN_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL__WILL_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL__imem_master_rready = RTL__near_mem$imem_master_rready ; 
  assign  RTL__dmem_master_awvalid = RTL__near_mem$dmem_master_awvalid ; 
  assign  RTL__dmem_master_awid = RTL__near_mem$dmem_master_awid ; 
  assign  RTL__dmem_master_awaddr = RTL__near_mem$dmem_master_awaddr ; 
  assign  RTL__dmem_master_awlen = RTL__near_mem$dmem_master_awlen ; 
  assign  RTL__dmem_master_awsize = RTL__near_mem$dmem_master_awsize ; 
  assign  RTL__dmem_master_awburst = RTL__near_mem$dmem_master_awburst ; 
  assign  RTL__dmem_master_awlock = RTL__near_mem$dmem_master_awlock ; 
  assign  RTL__dmem_master_awcache = RTL__near_mem$dmem_master_awcache ; 
  assign  RTL__dmem_master_awprot = RTL__near_mem$dmem_master_awprot ; 
  assign  RTL__dmem_master_awqos = RTL__near_mem$dmem_master_awqos ; 
  assign  RTL__dmem_master_awregion = RTL__near_mem$dmem_master_awregion ; 
  assign  RTL__CAN_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL__WILL_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL__dmem_master_wvalid = RTL__near_mem$dmem_master_wvalid ; 
  assign  RTL__dmem_master_wdata = RTL__near_mem$dmem_master_wdata ; 
  assign  RTL__dmem_master_wstrb = RTL__near_mem$dmem_master_wstrb ; 
  assign  RTL__dmem_master_wlast = RTL__near_mem$dmem_master_wlast ; 
  assign  RTL__CAN_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL__WILL_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL__CAN_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL__WILL_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL__dmem_master_bready = RTL__near_mem$dmem_master_bready ; 
  assign  RTL__dmem_master_arvalid = RTL__near_mem$dmem_master_arvalid ; 
  assign  RTL__dmem_master_arid = RTL__near_mem$dmem_master_arid ; 
  assign  RTL__dmem_master_araddr = RTL__near_mem$dmem_master_araddr ; 
  assign  RTL__dmem_master_arlen = RTL__near_mem$dmem_master_arlen ; 
  assign  RTL__dmem_master_arsize = RTL__near_mem$dmem_master_arsize ; 
  assign  RTL__dmem_master_arburst = RTL__near_mem$dmem_master_arburst ; 
  assign  RTL__dmem_master_arlock = RTL__near_mem$dmem_master_arlock ; 
  assign  RTL__dmem_master_arcache = RTL__near_mem$dmem_master_arcache ; 
  assign  RTL__dmem_master_arprot = RTL__near_mem$dmem_master_arprot ; 
  assign  RTL__dmem_master_arqos = RTL__near_mem$dmem_master_arqos ; 
  assign  RTL__dmem_master_arregion = RTL__near_mem$dmem_master_arregion ; 
  assign  RTL__CAN_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL__WILL_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL__CAN_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL__WILL_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL__dmem_master_rready = RTL__near_mem$dmem_master_rready ; 
  assign  RTL__CAN_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL__WILL_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL__CAN_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL__WILL_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL__CAN_FIRE_software_interrupt_req =1'd1; 
  assign  RTL__WILL_FIRE_software_interrupt_req =1'd1; 
  assign  RTL__CAN_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL__WILL_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL__CAN_FIRE_nmi_req =1'd1; 
  assign  RTL__WILL_FIRE_nmi_req =1'd1; 
  assign  RTL__RDY_set_verbosity =1'd1; 
  assign  RTL__CAN_FIRE_set_verbosity =1'd1; 
  assign  RTL__WILL_FIRE_set_verbosity = RTL__EN_set_verbosity ;  
    wire RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__rg_nmi;
    wire RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__rg_state;
    wire RTL__csr_regfile__CLK;
    wire RTL__csr_regfile__RST_N;
    wire RTL__csr_regfile__EN_server_reset_request_put;
    wire RTL__csr_regfile__RDY_server_reset_request_put;
    wire RTL__csr_regfile__EN_server_reset_response_get;
    wire RTL__csr_regfile__RDY_server_reset_response_get;
    wire[11:0] RTL__csr_regfile__read_csr_csr_addr;
    wire[32:0] RTL__csr_regfile__read_csr;
    wire[11:0] RTL__csr_regfile__read_csr_port2_csr_addr;
    wire[32:0] RTL__csr_regfile__read_csr_port2;
    wire[11:0] RTL__csr_regfile__mav_read_csr_csr_addr;
    wire RTL__csr_regfile__EN_mav_read_csr;
    wire[32:0] RTL__csr_regfile__mav_read_csr;
    wire[11:0] RTL__csr_regfile__mav_csr_write_csr_addr;
    wire[31:0] RTL__csr_regfile__mav_csr_write_word;
    wire RTL__csr_regfile__EN_mav_csr_write;
    wire[31:0] RTL__csr_regfile__mav_csr_write;
    wire[27:0] RTL__csr_regfile__read_misa;
    wire[31:0] RTL__csr_regfile__read_mstatus;
    wire[31:0] RTL__csr_regfile__read_ustatus;
    wire[31:0] RTL__csr_regfile__read_satp;
    wire[1:0] RTL__csr_regfile__csr_trap_actions_from_priv;
    wire[31:0] RTL__csr_regfile__csr_trap_actions_pc;
    wire RTL__csr_regfile__csr_trap_actions_nmi;
    wire RTL__csr_regfile__csr_trap_actions_interrupt;
    wire[3:0] RTL__csr_regfile__csr_trap_actions_exc_code;
    wire[31:0] RTL__csr_regfile__csr_trap_actions_xtval;
    wire RTL__csr_regfile__EN_csr_trap_actions;
    wire[97:0] RTL__csr_regfile__csr_trap_actions;
    wire RTL__csr_regfile__RDY_csr_trap_actions;
    wire[1:0] RTL__csr_regfile__csr_ret_actions_from_priv;
    wire RTL__csr_regfile__EN_csr_ret_actions;
    wire[65:0] RTL__csr_regfile__csr_ret_actions;
    wire RTL__csr_regfile__RDY_csr_ret_actions;
    wire[63:0] RTL__csr_regfile__read_csr_minstret;
    wire RTL__csr_regfile__EN_csr_minstret_incr;
    wire[63:0] RTL__csr_regfile__read_csr_mcycle;
    wire[63:0] RTL__csr_regfile__read_csr_mtime;
    wire[1:0] RTL__csr_regfile__access_permitted_1_priv;
    wire[11:0] RTL__csr_regfile__access_permitted_1_csr_addr;
    wire RTL__csr_regfile__access_permitted_1_read_not_write;
    wire RTL__csr_regfile__access_permitted_1;
    wire[1:0] RTL__csr_regfile__access_permitted_2_priv;
    wire[11:0] RTL__csr_regfile__access_permitted_2_csr_addr;
    wire RTL__csr_regfile__access_permitted_2_read_not_write;
    wire RTL__csr_regfile__access_permitted_2;
    wire[1:0] RTL__csr_regfile__csr_counter_read_fault_priv;
    wire[11:0] RTL__csr_regfile__csr_counter_read_fault_csr_addr;
    wire RTL__csr_regfile__csr_counter_read_fault;
    wire[31:0] RTL__csr_regfile__csr_mip_read;
    wire RTL__csr_regfile__m_external_interrupt_req_set_not_clear;
    wire RTL__csr_regfile__s_external_interrupt_req_set_not_clear;
    wire RTL__csr_regfile__timer_interrupt_req_set_not_clear;
    wire RTL__csr_regfile__software_interrupt_req_set_not_clear;
    wire[1:0] RTL__csr_regfile__interrupt_pending_cur_priv;
    wire[4:0] RTL__csr_regfile__interrupt_pending;
    wire RTL__csr_regfile__wfi_resume;
    wire RTL__csr_regfile__nmi_req_set_not_clear;
    wire RTL__csr_regfile__nmi_pending;
    wire RTL__csr_regfile__EN_debug;
    wire RTL__csr_regfile__RDY_debug;

    wire[97:0] RTL__csr_regfile__csr_trap_actions ; 
    wire[65:0] RTL__csr_regfile__csr_ret_actions ; 
    wire[63:0] RTL__csr_regfile__read_csr_mcycle , RTL__csr_regfile__read_csr_minstret , RTL__csr_regfile__read_csr_mtime ; 
    wire[32:0] RTL__csr_regfile__mav_read_csr , RTL__csr_regfile__read_csr , RTL__csr_regfile__read_csr_port2 ; 
    wire[31:0] RTL__csr_regfile__csr_mip_read , RTL__csr_regfile__mav_csr_write , RTL__csr_regfile__read_mstatus , RTL__csr_regfile__read_satp , RTL__csr_regfile__read_ustatus ; 
    wire[27:0] RTL__csr_regfile__read_misa ; 
    wire[4:0] RTL__csr_regfile__interrupt_pending ; 
    wire RTL__csr_regfile__RDY_csr_ret_actions , RTL__csr_regfile__RDY_csr_trap_actions , RTL__csr_regfile__RDY_debug , RTL__csr_regfile__RDY_server_reset_request_put , RTL__csr_regfile__RDY_server_reset_response_get , RTL__csr_regfile__access_permitted_1 , RTL__csr_regfile__access_permitted_2 , RTL__csr_regfile__csr_counter_read_fault , RTL__csr_regfile__nmi_pending , RTL__csr_regfile__wfi_resume ; reg[3:0] RTL__csr_regfile__cfg_verbosity ; 
    wire[3:0] RTL__csr_regfile__cfg_verbosity$D_IN ; 
    wire RTL__csr_regfile__cfg_verbosity$EN ; reg[31:0] RTL__csr_regfile__csr_mstatus_rg_mstatus ; reg[31:0] RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN ; 
    wire RTL__csr_regfile__csr_mstatus_rg_mstatus$EN ; reg[31:0] RTL__csr_regfile__rg_dcsr ; 
    wire[31:0] RTL__csr_regfile__rg_dcsr$D_IN ; 
    wire RTL__csr_regfile__rg_dcsr$EN ; reg[31:0] RTL__csr_regfile__rg_dpc ; 
    wire[31:0] RTL__csr_regfile__rg_dpc$D_IN ; 
    wire RTL__csr_regfile__rg_dpc$EN ; reg[31:0] RTL__csr_regfile__rg_dscratch0 ; 
    wire[31:0] RTL__csr_regfile__rg_dscratch0$D_IN ; 
    wire RTL__csr_regfile__rg_dscratch0$EN ; reg[31:0] RTL__csr_regfile__rg_dscratch1 ; 
    wire[31:0] RTL__csr_regfile__rg_dscratch1$D_IN ; 
    wire RTL__csr_regfile__rg_dscratch1$EN ; reg[4:0] RTL__csr_regfile__rg_mcause ; reg[4:0] RTL__csr_regfile__rg_mcause$D_IN ; 
    wire RTL__csr_regfile__rg_mcause$EN ; reg[2:0] RTL__csr_regfile__rg_mcounteren ; 
    wire[2:0] RTL__csr_regfile__rg_mcounteren$D_IN ; 
    wire RTL__csr_regfile__rg_mcounteren$EN ; reg[63:0] RTL__csr_regfile__rg_mcycle ; 
    wire[63:0] RTL__csr_regfile__rg_mcycle$D_IN ; 
    wire RTL__csr_regfile__rg_mcycle$EN ; reg[31:0] RTL__csr_regfile__rg_mepc ; 
    wire[31:0] RTL__csr_regfile__rg_mepc$D_IN ; 
    wire RTL__csr_regfile__rg_mepc$EN ; reg[63:0] RTL__csr_regfile__rg_minstret ; 
    wire[63:0] RTL__csr_regfile__rg_minstret$D_IN ; 
    wire RTL__csr_regfile__rg_minstret$EN ; reg[31:0] RTL__csr_regfile__rg_mscratch ; 
    wire[31:0] RTL__csr_regfile__rg_mscratch$D_IN ; 
    wire RTL__csr_regfile__rg_mscratch$EN ; reg[31:0] RTL__csr_regfile__rg_mtval ; 
    wire[31:0] RTL__csr_regfile__rg_mtval$D_IN ; 
    wire RTL__csr_regfile__rg_mtval$EN ; reg[30:0] RTL__csr_regfile__rg_mtvec ; 
    wire[30:0] RTL__csr_regfile__rg_mtvec$D_IN ; 
    wire RTL__csr_regfile__rg_mtvec$EN ; 
    reg RTL__csr_regfile__rg_nmi ; 
    wire RTL__csr_regfile__rg_nmi$D_IN , RTL__csr_regfile__rg_nmi$EN ; reg[31:0] RTL__csr_regfile__rg_nmi_vector ; 
    wire[31:0] RTL__csr_regfile__rg_nmi_vector$D_IN ; 
    wire RTL__csr_regfile__rg_nmi_vector$EN ; 
    reg RTL__csr_regfile__rg_state ; 
    wire RTL__csr_regfile__rg_state$D_IN , RTL__csr_regfile__rg_state$EN ; reg[31:0] RTL__csr_regfile__rg_tdata1 ; 
    wire[31:0] RTL__csr_regfile__rg_tdata1$D_IN ; 
    wire RTL__csr_regfile__rg_tdata1$EN ; reg[31:0] RTL__csr_regfile__rg_tdata2 ; 
    wire[31:0] RTL__csr_regfile__rg_tdata2$D_IN ; 
    wire RTL__csr_regfile__rg_tdata2$EN ; reg[31:0] RTL__csr_regfile__rg_tdata3 ; 
    wire[31:0] RTL__csr_regfile__rg_tdata3$D_IN ; 
    wire RTL__csr_regfile__rg_tdata3$EN ; reg[31:0] RTL__csr_regfile__rg_tselect ; 
    wire[31:0] RTL__csr_regfile__rg_tselect$D_IN ; 
    wire RTL__csr_regfile__rg_tselect$EN ; 
    wire[31:0] RTL__csr_regfile__csr_mie$fav_write , RTL__csr_regfile__csr_mie$fav_write_wordxl , RTL__csr_regfile__csr_mie$fv_read ; 
    wire[27:0] RTL__csr_regfile__csr_mie$fav_write_misa ; 
    wire RTL__csr_regfile__csr_mie$EN_fav_write , RTL__csr_regfile__csr_mie$EN_reset ; 
    wire[31:0] RTL__csr_regfile__csr_mip$fav_write , RTL__csr_regfile__csr_mip$fav_write_wordxl , RTL__csr_regfile__csr_mip$fv_read ; 
    wire[27:0] RTL__csr_regfile__csr_mip$fav_write_misa ; 
    wire RTL__csr_regfile__csr_mip$EN_fav_write , RTL__csr_regfile__csr_mip$EN_reset , RTL__csr_regfile__csr_mip$m_external_interrupt_req_req , RTL__csr_regfile__csr_mip$s_external_interrupt_req_req , RTL__csr_regfile__csr_mip$software_interrupt_req_req , RTL__csr_regfile__csr_mip$timer_interrupt_req_req ; 
    wire RTL__csr_regfile__f_reset_rsps$CLR , RTL__csr_regfile__f_reset_rsps$DEQ , RTL__csr_regfile__f_reset_rsps$EMPTY_N , RTL__csr_regfile__f_reset_rsps$ENQ , RTL__csr_regfile__f_reset_rsps$FULL_N ; 
    wire[63:0] RTL__csr_regfile__soc_map$m_is_IO_addr_addr , RTL__csr_regfile__soc_map$m_is_mem_addr_addr , RTL__csr_regfile__soc_map$m_is_near_mem_IO_addr_addr , RTL__csr_regfile__soc_map$m_mtvec_reset_value , RTL__csr_regfile__soc_map$m_nmivec_reset_value ; 
    wire RTL__csr_regfile__CAN_FIRE_RL_rl_mcycle_incr , RTL__csr_regfile__CAN_FIRE_RL_rl_reset_start , RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_csrrx , RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_incr , RTL__csr_regfile__CAN_FIRE_csr_minstret_incr , RTL__csr_regfile__CAN_FIRE_csr_ret_actions , RTL__csr_regfile__CAN_FIRE_csr_trap_actions , RTL__csr_regfile__CAN_FIRE_debug , RTL__csr_regfile__CAN_FIRE_m_external_interrupt_req , RTL__csr_regfile__CAN_FIRE_mav_csr_write , RTL__csr_regfile__CAN_FIRE_mav_read_csr , RTL__csr_regfile__CAN_FIRE_nmi_req , RTL__csr_regfile__CAN_FIRE_s_external_interrupt_req , RTL__csr_regfile__CAN_FIRE_server_reset_request_put , RTL__csr_regfile__CAN_FIRE_server_reset_response_get , RTL__csr_regfile__CAN_FIRE_software_interrupt_req , RTL__csr_regfile__CAN_FIRE_timer_interrupt_req , RTL__csr_regfile__WILL_FIRE_RL_rl_mcycle_incr , RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start , RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_csrrx , RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_incr , RTL__csr_regfile__WILL_FIRE_csr_minstret_incr , RTL__csr_regfile__WILL_FIRE_csr_ret_actions , RTL__csr_regfile__WILL_FIRE_csr_trap_actions , RTL__csr_regfile__WILL_FIRE_debug , RTL__csr_regfile__WILL_FIRE_m_external_interrupt_req , RTL__csr_regfile__WILL_FIRE_mav_csr_write , RTL__csr_regfile__WILL_FIRE_mav_read_csr , RTL__csr_regfile__WILL_FIRE_nmi_req , RTL__csr_regfile__WILL_FIRE_s_external_interrupt_req , RTL__csr_regfile__WILL_FIRE_server_reset_request_put , RTL__csr_regfile__WILL_FIRE_server_reset_response_get , RTL__csr_regfile__WILL_FIRE_software_interrupt_req , RTL__csr_regfile__WILL_FIRE_timer_interrupt_req ; 
    wire[63:0] RTL__csr_regfile__MUX_rg_minstret$write_1__VAL_1 , RTL__csr_regfile__MUX_rg_minstret$write_1__VAL_2 , RTL__csr_regfile__MUX_rw_minstret$wset_1__VAL_1 ; 
    wire[31:0] RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__VAL_3 ; 
    wire[30:0] RTL__csr_regfile__MUX_rg_mtvec$write_1__VAL_1 , RTL__csr_regfile__MUX_rg_mtvec$write_1__VAL_2 ; 
    wire[4:0] RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_2 , RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_3 ; 
    wire RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__SEL_2 , RTL__csr_regfile__MUX_rg_mcause$write_1__SEL_2 , RTL__csr_regfile__MUX_rg_mcounteren$write_1__SEL_1 , RTL__csr_regfile__MUX_rg_mepc$write_1__SEL_1 , RTL__csr_regfile__MUX_rg_mtval$write_1__SEL_1 , RTL__csr_regfile__MUX_rg_mtvec$write_1__SEL_1 , RTL__csr_regfile__MUX_rg_state$write_1__SEL_2 , RTL__csr_regfile__MUX_rg_tdata1$write_1__SEL_1 , RTL__csr_regfile__MUX_rw_minstret$wset_1__SEL_1 ; reg[31:0] RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769 , RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574 , RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220 , RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397 ; 
    wire[63:0] RTL__csr_regfile__x__h5174 , RTL__csr_regfile__x__h5282 ; 
    wire[33:0] RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1068 ; 
    wire[31:0] RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 , RTL__csr_regfile___theResult___fst__h8211 , RTL__csr_regfile___theResult___fst__h8412 , RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 , RTL__csr_regfile__exc_pc___1__h7296 , RTL__csr_regfile__exc_pc__h7032 , RTL__csr_regfile__exc_pc__h7243 , RTL__csr_regfile__mask__h8232 , RTL__csr_regfile__mask__h8249 , RTL__csr_regfile__result__h4701 , RTL__csr_regfile__result__h5357 , RTL__csr_regfile__v__h4509 , RTL__csr_regfile__v__h4571 , RTL__csr_regfile__v__h4742 , RTL__csr_regfile__val__h8250 , RTL__csr_regfile__vector_offset__h7244 , RTL__csr_regfile__wordxl1__h4038 , RTL__csr_regfile__x__h5843 , RTL__csr_regfile__x__h8067 , RTL__csr_regfile__x__h8068 , RTL__csr_regfile__x__h8085 , RTL__csr_regfile__x__h8231 , RTL__csr_regfile__x__h8244 , RTL__csr_regfile__x__h8261 , RTL__csr_regfile__y__h8245 , RTL__csr_regfile__y__h8262 ; 
    wire[22:0] RTL__csr_regfile__fixed_up_val_23__h4079 , RTL__csr_regfile__fixed_up_val_23__h6471 , RTL__csr_regfile__fixed_up_val_23__h8130 ; 
    wire[5:0] RTL__csr_regfile__ie_from_x__h8195 , RTL__csr_regfile__pie_from_x__h8196 ; 
    wire[3:0] RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1370 , RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1372 , RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1374 , RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1376 , RTL__csr_regfile__exc_code__h7909 ; 
    wire[1:0] RTL__csr_regfile__mpp__h7337 , RTL__csr_regfile__to_y__h8411 ; 
    wire RTL__csr_regfile__NOT_access_permitted_1_csr_addr_ULT_0xC03_069__ETC___d1155 , RTL__csr_regfile__NOT_access_permitted_2_csr_addr_ULT_0xC03_160__ETC___d1245 , RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1364 , RTL__csr_regfile__NOT_csr_trap_actions_nmi_97_AND_csr_trap_actio_ETC___d974 , RTL__csr_regfile__NOT_mav_csr_write_csr_addr_ULT_0xB03_77_35_AND_ETC___d746 , RTL__csr_regfile__b__h8248 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1288 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1293 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1298 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1303 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1308 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1313 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1318 , RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1323 , RTL__csr_regfile__csr_trap_actions_nmi_OR_NOT_csr_trap_actions_i_ETC___d1025 , RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0x33F___d586 , RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB1F___d578 , RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB9F___d582 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323_85_OR_NOT_mav_ETC___d728 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323___d585 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d642 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d730 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03___d577 , RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB83___d581 ; 
  assign  RTL__csr_regfile__RDY_server_reset_request_put = RTL__csr_regfile__f_reset_rsps$FULL_N ; 
  assign  RTL__csr_regfile__CAN_FIRE_server_reset_request_put = RTL__csr_regfile__f_reset_rsps$FULL_N ; 
  assign  RTL__csr_regfile__WILL_FIRE_server_reset_request_put = RTL__csr_regfile__EN_server_reset_request_put ; 
  assign  RTL__csr_regfile__RDY_server_reset_response_get = RTL__csr_regfile__rg_state && RTL__csr_regfile__f_reset_rsps$EMPTY_N ; 
  assign  RTL__csr_regfile__CAN_FIRE_server_reset_response_get = RTL__csr_regfile__rg_state && RTL__csr_regfile__f_reset_rsps$EMPTY_N ; 
  assign  RTL__csr_regfile__WILL_FIRE_server_reset_response_get = RTL__csr_regfile__EN_server_reset_response_get ; 
  assign  RTL__csr_regfile__read_csr ={ RTL__csr_regfile__read_csr_csr_addr >=12'hC03&& RTL__csr_regfile__read_csr_csr_addr <=12'hC1F|| RTL__csr_regfile__read_csr_csr_addr >=12'hC83&& RTL__csr_regfile__read_csr_csr_addr <=12'hC9F|| RTL__csr_regfile__read_csr_csr_addr >=12'hB03&& RTL__csr_regfile__read_csr_csr_addr <=12'hB1F|| RTL__csr_regfile__read_csr_csr_addr >=12'hB83&& RTL__csr_regfile__read_csr_csr_addr <=12'hB9F|| RTL__csr_regfile__read_csr_csr_addr >=12'h323&& RTL__csr_regfile__read_csr_csr_addr <=12'h33F|| RTL__csr_regfile__read_csr_csr_addr ==12'hC00|| RTL__csr_regfile__read_csr_csr_addr ==12'hC02|| RTL__csr_regfile__read_csr_csr_addr ==12'hC80|| RTL__csr_regfile__read_csr_csr_addr ==12'hC82|| RTL__csr_regfile__read_csr_csr_addr ==12'hF11|| RTL__csr_regfile__read_csr_csr_addr ==12'hF12|| RTL__csr_regfile__read_csr_csr_addr ==12'hF13|| RTL__csr_regfile__read_csr_csr_addr ==12'hF14|| RTL__csr_regfile__read_csr_csr_addr ==12'h300|| RTL__csr_regfile__read_csr_csr_addr ==12'h301|| RTL__csr_regfile__read_csr_csr_addr ==12'h304|| RTL__csr_regfile__read_csr_csr_addr ==12'h305|| RTL__csr_regfile__read_csr_csr_addr ==12'h306|| RTL__csr_regfile__read_csr_csr_addr ==12'h340|| RTL__csr_regfile__read_csr_csr_addr ==12'h341|| RTL__csr_regfile__read_csr_csr_addr ==12'h342|| RTL__csr_regfile__read_csr_csr_addr ==12'h343|| RTL__csr_regfile__read_csr_csr_addr ==12'h344|| RTL__csr_regfile__read_csr_csr_addr ==12'hB00|| RTL__csr_regfile__read_csr_csr_addr ==12'hB02|| RTL__csr_regfile__read_csr_csr_addr ==12'hB80|| RTL__csr_regfile__read_csr_csr_addr ==12'hB82|| RTL__csr_regfile__read_csr_csr_addr ==12'h7A0|| RTL__csr_regfile__read_csr_csr_addr ==12'h7A1|| RTL__csr_regfile__read_csr_csr_addr ==12'h7A2|| RTL__csr_regfile__read_csr_csr_addr ==12'h7A3,( RTL__csr_regfile__read_csr_csr_addr >=12'hC03&& RTL__csr_regfile__read_csr_csr_addr <=12'hC1F|| RTL__csr_regfile__read_csr_csr_addr >=12'hC83&& RTL__csr_regfile__read_csr_csr_addr <=12'hC9F|| RTL__csr_regfile__read_csr_csr_addr >=12'hB03&& RTL__csr_regfile__read_csr_csr_addr <=12'hB1F|| RTL__csr_regfile__read_csr_csr_addr >=12'hB83&& RTL__csr_regfile__read_csr_csr_addr <=12'hB9F|| RTL__csr_regfile__read_csr_csr_addr >=12'h323&& RTL__csr_regfile__read_csr_csr_addr <=12'h33F) ? 32'd0: RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220 }; 
  assign  RTL__csr_regfile__read_csr_port2 ={ RTL__csr_regfile__read_csr_port2_csr_addr >=12'hC03&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hC1F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'hC83&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hC9F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'hB03&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hB1F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'hB83&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hB9F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'h323&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'h33F|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hC00|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hC02|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hC80|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hC82|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hF11|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hF12|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hF13|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hF14|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h300|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h301|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h304|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h305|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h306|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h340|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h341|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h342|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h343|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h344|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hB00|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hB02|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hB80|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'hB82|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h7A0|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h7A1|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h7A2|| RTL__csr_regfile__read_csr_port2_csr_addr ==12'h7A3,( RTL__csr_regfile__read_csr_port2_csr_addr >=12'hC03&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hC1F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'hC83&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hC9F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'hB03&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hB1F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'hB83&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'hB9F|| RTL__csr_regfile__read_csr_port2_csr_addr >=12'h323&& RTL__csr_regfile__read_csr_port2_csr_addr <=12'h33F) ? 32'd0: RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397 }; 
  assign  RTL__csr_regfile__mav_read_csr ={ RTL__csr_regfile__mav_read_csr_csr_addr >=12'hC03&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hC1F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'hC83&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hC9F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'hB03&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hB1F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'hB83&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hB9F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'h323&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'h33F|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hC00|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hC02|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hC80|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hC82|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hF11|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hF12|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hF13|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hF14|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h300|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h301|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h304|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h305|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h306|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h340|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h341|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h342|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h343|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h344|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hB00|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hB02|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hB80|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'hB82|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h7A0|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h7A1|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h7A2|| RTL__csr_regfile__mav_read_csr_csr_addr ==12'h7A3,( RTL__csr_regfile__mav_read_csr_csr_addr >=12'hC03&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hC1F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'hC83&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hC9F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'hB03&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hB1F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'hB83&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'hB9F|| RTL__csr_regfile__mav_read_csr_csr_addr >=12'h323&& RTL__csr_regfile__mav_read_csr_csr_addr <=12'h33F) ? 32'd0: RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574 }; 
  assign  RTL__csr_regfile__CAN_FIRE_mav_read_csr =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_mav_read_csr = RTL__csr_regfile__EN_mav_read_csr ; 
  assign  RTL__csr_regfile__mav_csr_write = RTL__csr_regfile__NOT_mav_csr_write_csr_addr_ULT_0xB03_77_35_AND_ETC___d746  ? 32'd0: RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769 ; 
  assign  RTL__csr_regfile__CAN_FIRE_mav_csr_write =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_mav_csr_write = RTL__csr_regfile__EN_mav_csr_write ; 
  assign  RTL__csr_regfile__read_misa =28'd68157696; 
  assign  RTL__csr_regfile__read_mstatus = RTL__csr_regfile__csr_mstatus_rg_mstatus ; 
  assign  RTL__csr_regfile__read_ustatus ={27'd0, RTL__csr_regfile__csr_mstatus_rg_mstatus [4],3'd0, RTL__csr_regfile__csr_mstatus_rg_mstatus [0]}; 
  assign  RTL__csr_regfile__read_satp =32'hAAAAAAAA; 
  assign  RTL__csr_regfile__csr_trap_actions ={ RTL__csr_regfile__x__h5843 , RTL__csr_regfile__x__h8067 , RTL__csr_regfile__x__h8068 ,2'b11}; 
  assign  RTL__csr_regfile__RDY_csr_trap_actions =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_csr_trap_actions =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_csr_trap_actions = RTL__csr_regfile__EN_csr_trap_actions ; 
  assign  RTL__csr_regfile__csr_ret_actions ={ RTL__csr_regfile__x__h8085 , RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1068 }; 
  assign  RTL__csr_regfile__RDY_csr_ret_actions =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_csr_ret_actions =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_csr_ret_actions = RTL__csr_regfile__EN_csr_ret_actions ; 
  assign  RTL__csr_regfile__read_csr_minstret = RTL__csr_regfile__rg_minstret ; 
  assign  RTL__csr_regfile__CAN_FIRE_csr_minstret_incr =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_csr_minstret_incr = RTL__csr_regfile__EN_csr_minstret_incr ; 
  assign  RTL__csr_regfile__read_csr_mcycle = RTL__csr_regfile__rg_mcycle ; 
  assign  RTL__csr_regfile__read_csr_mtime = RTL__csr_regfile__rg_mcycle ; 
  assign  RTL__csr_regfile__access_permitted_1 = RTL__csr_regfile__NOT_access_permitted_1_csr_addr_ULT_0xC03_069__ETC___d1155 &&( RTL__csr_regfile__access_permitted_1_read_not_write || RTL__csr_regfile__access_permitted_1_csr_addr [11:10]!=2'b11); 
  assign  RTL__csr_regfile__access_permitted_2 = RTL__csr_regfile__NOT_access_permitted_2_csr_addr_ULT_0xC03_160__ETC___d1245 &&( RTL__csr_regfile__access_permitted_2_read_not_write || RTL__csr_regfile__access_permitted_2_csr_addr [11:10]!=2'b11); 
  assign  RTL__csr_regfile__csr_counter_read_fault =( RTL__csr_regfile__csr_counter_read_fault_priv ==2'b01|| RTL__csr_regfile__csr_counter_read_fault_priv ==2'b0)&&( RTL__csr_regfile__csr_counter_read_fault_csr_addr ==12'hC00&&! RTL__csr_regfile__rg_mcounteren [0]|| RTL__csr_regfile__csr_counter_read_fault_csr_addr ==12'hC01&&! RTL__csr_regfile__rg_mcounteren [1]|| RTL__csr_regfile__csr_counter_read_fault_csr_addr ==12'hC02&&! RTL__csr_regfile__rg_mcounteren [2]|| RTL__csr_regfile__csr_counter_read_fault_csr_addr >=12'hC03&& RTL__csr_regfile__csr_counter_read_fault_csr_addr <=12'hC1F|| RTL__csr_regfile__csr_counter_read_fault_csr_addr >=12'hC83&& RTL__csr_regfile__csr_counter_read_fault_csr_addr <=12'hC9F); 
  assign  RTL__csr_regfile__csr_mip_read = RTL__csr_regfile__csr_mip$fv_read ; 
  assign  RTL__csr_regfile__CAN_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_software_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_software_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__interrupt_pending ={ RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1323 , RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1364  ? 4'd4: RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1376 }; 
  assign  RTL__csr_regfile__wfi_resume =( RTL__csr_regfile__csr_mip$fv_read & RTL__csr_regfile__csr_mie$fv_read )!=32'd0; 
  assign  RTL__csr_regfile__CAN_FIRE_nmi_req =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_nmi_req =1'd1; 
  assign  RTL__csr_regfile__nmi_pending = RTL__csr_regfile__rg_nmi ; 
  assign  RTL__csr_regfile__RDY_debug =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_debug =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_debug = RTL__csr_regfile__EN_debug ;  
    wire RTL__csr_regfile__csr_mie__CLK;
    wire RTL__csr_regfile__csr_mie__RST_N;
    wire RTL__csr_regfile__csr_mie__EN_reset;
    wire[31:0] RTL__csr_regfile__csr_mie__fv_read;
    wire[27:0] RTL__csr_regfile__csr_mie__fav_write_misa;
    wire[31:0] RTL__csr_regfile__csr_mie__fav_write_wordxl;
    wire RTL__csr_regfile__csr_mie__EN_fav_write;
    wire[31:0] RTL__csr_regfile__csr_mie__fav_write;

    wire[31:0] RTL__csr_regfile__csr_mie__fav_write , RTL__csr_regfile__csr_mie__fv_read ; reg[11:0] RTL__csr_regfile__csr_mie__rg_mie ; 
    wire[11:0] RTL__csr_regfile__csr_mie__rg_mie$D_IN ; 
    wire RTL__csr_regfile__csr_mie__rg_mie$EN ; 
    wire RTL__csr_regfile__csr_mie__CAN_FIRE_fav_write , RTL__csr_regfile__csr_mie__CAN_FIRE_reset , RTL__csr_regfile__csr_mie__WILL_FIRE_fav_write , RTL__csr_regfile__csr_mie__WILL_FIRE_reset ; 
    wire[11:0] RTL__csr_regfile__csr_mie__mie__h88 ; 
    wire RTL__csr_regfile__csr_mie__seie__h119 , RTL__csr_regfile__csr_mie__ssie__h113 , RTL__csr_regfile__csr_mie__stie__h116 , RTL__csr_regfile__csr_mie__ueie__h118 , RTL__csr_regfile__csr_mie__usie__h112 , RTL__csr_regfile__csr_mie__utie__h115 ; 
  assign  RTL__csr_regfile__csr_mie__CAN_FIRE_reset =1'd1; 
  assign  RTL__csr_regfile__csr_mie__WILL_FIRE_reset = RTL__csr_regfile__csr_mie__EN_reset ; 
  assign  RTL__csr_regfile__csr_mie__fv_read ={20'd0, RTL__csr_regfile__csr_mie__rg_mie }; 
  assign  RTL__csr_regfile__csr_mie__fav_write ={20'd0, RTL__csr_regfile__csr_mie__mie__h88 }; 
  assign  RTL__csr_regfile__csr_mie__CAN_FIRE_fav_write =1'd1; 
  assign  RTL__csr_regfile__csr_mie__WILL_FIRE_fav_write = RTL__csr_regfile__csr_mie__EN_fav_write ; 
  assign  RTL__csr_regfile__csr_mie__rg_mie$D_IN = RTL__csr_regfile__csr_mie__EN_fav_write  ?  RTL__csr_regfile__csr_mie__mie__h88 :12'd0; 
  assign  RTL__csr_regfile__csr_mie__rg_mie$EN = RTL__csr_regfile__csr_mie__EN_fav_write || RTL__csr_regfile__csr_mie__EN_reset ; 
  assign  RTL__csr_regfile__csr_mie__mie__h88 ={ RTL__csr_regfile__csr_mie__fav_write_wordxl [11],1'b0, RTL__csr_regfile__csr_mie__seie__h119 , RTL__csr_regfile__csr_mie__ueie__h118 , RTL__csr_regfile__csr_mie__fav_write_wordxl [7],1'b0, RTL__csr_regfile__csr_mie__stie__h116 , RTL__csr_regfile__csr_mie__utie__h115 , RTL__csr_regfile__csr_mie__fav_write_wordxl [3],1'b0, RTL__csr_regfile__csr_mie__ssie__h113 , RTL__csr_regfile__csr_mie__usie__h112 }; 
  assign  RTL__csr_regfile__csr_mie__seie__h119 = RTL__csr_regfile__csr_mie__fav_write_misa [18]&& RTL__csr_regfile__csr_mie__fav_write_wordxl [9]; 
  assign  RTL__csr_regfile__csr_mie__ssie__h113 = RTL__csr_regfile__csr_mie__fav_write_misa [18]&& RTL__csr_regfile__csr_mie__fav_write_wordxl [1]; 
  assign  RTL__csr_regfile__csr_mie__stie__h116 = RTL__csr_regfile__csr_mie__fav_write_misa [18]&& RTL__csr_regfile__csr_mie__fav_write_wordxl [5]; 
  assign  RTL__csr_regfile__csr_mie__ueie__h118 = RTL__csr_regfile__csr_mie__fav_write_misa [13]&& RTL__csr_regfile__csr_mie__fav_write_wordxl [8]; 
  assign  RTL__csr_regfile__csr_mie__usie__h112 = RTL__csr_regfile__csr_mie__fav_write_misa [13]&& RTL__csr_regfile__csr_mie__fav_write_wordxl [0]; 
  assign  RTL__csr_regfile__csr_mie__utie__h115 = RTL__csr_regfile__csr_mie__fav_write_misa [13]&& RTL__csr_regfile__csr_mie__fav_write_wordxl [4]; 
  always @( posedge  RTL__csr_regfile__csr_mie__CLK )
         begin 
             if ( RTL__csr_regfile__csr_mie__RST_N ==1'b0)
                 begin  
                     RTL__csr_regfile__csr_mie__rg_mie  <=12'd0;
                 end 
              else 
                 begin 
                     if ( RTL__csr_regfile__csr_mie__rg_mie$EN ) 
                         RTL__csr_regfile__csr_mie__rg_mie  <= RTL__csr_regfile__csr_mie__rg_mie$D_IN ;
                 end 
         end
 
    assign RTL__csr_regfile__csr_mie__CLK = RTL__csr_regfile__CLK;
    assign RTL__csr_regfile__csr_mie__RST_N = RTL__csr_regfile__RST_N;
    assign RTL__csr_regfile__csr_mie__EN_reset = RTL__csr_regfile__csr_mie$EN_reset;
    assign RTL__csr_regfile__csr_mie$fv_read = RTL__csr_regfile__csr_mie__fv_read;
    assign RTL__csr_regfile__csr_mie__fav_write_misa = RTL__csr_regfile__csr_mie$fav_write_misa;
    assign RTL__csr_regfile__csr_mie__fav_write_wordxl = RTL__csr_regfile__csr_mie$fav_write_wordxl;
    assign RTL__csr_regfile__csr_mie__EN_fav_write = RTL__csr_regfile__csr_mie$EN_fav_write;
    assign RTL__csr_regfile__csr_mie$fav_write = RTL__csr_regfile__csr_mie__fav_write;
      
    wire RTL__csr_regfile__csr_mip__CLK;
    wire RTL__csr_regfile__csr_mip__RST_N;
    wire RTL__csr_regfile__csr_mip__EN_reset;
    wire[31:0] RTL__csr_regfile__csr_mip__fv_read;
    wire[27:0] RTL__csr_regfile__csr_mip__fav_write_misa;
    wire[31:0] RTL__csr_regfile__csr_mip__fav_write_wordxl;
    wire RTL__csr_regfile__csr_mip__EN_fav_write;
    wire[31:0] RTL__csr_regfile__csr_mip__fav_write;
    wire RTL__csr_regfile__csr_mip__m_external_interrupt_req_req;
    wire RTL__csr_regfile__csr_mip__s_external_interrupt_req_req;
    wire RTL__csr_regfile__csr_mip__software_interrupt_req_req;
    wire RTL__csr_regfile__csr_mip__timer_interrupt_req_req;

    wire[31:0] RTL__csr_regfile__csr_mip__fav_write , RTL__csr_regfile__csr_mip__fv_read ; 
    reg RTL__csr_regfile__csr_mip__rg_meip ; 
    wire RTL__csr_regfile__csr_mip__rg_meip$D_IN , RTL__csr_regfile__csr_mip__rg_meip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_msip ; 
    wire RTL__csr_regfile__csr_mip__rg_msip$D_IN , RTL__csr_regfile__csr_mip__rg_msip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_mtip ; 
    wire RTL__csr_regfile__csr_mip__rg_mtip$D_IN , RTL__csr_regfile__csr_mip__rg_mtip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_seip ; 
    wire RTL__csr_regfile__csr_mip__rg_seip$D_IN , RTL__csr_regfile__csr_mip__rg_seip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_ssip ; 
    wire RTL__csr_regfile__csr_mip__rg_ssip$D_IN , RTL__csr_regfile__csr_mip__rg_ssip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_stip ; 
    wire RTL__csr_regfile__csr_mip__rg_stip$D_IN , RTL__csr_regfile__csr_mip__rg_stip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_ueip ; 
    wire RTL__csr_regfile__csr_mip__rg_ueip$D_IN , RTL__csr_regfile__csr_mip__rg_ueip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_usip ; 
    wire RTL__csr_regfile__csr_mip__rg_usip$D_IN , RTL__csr_regfile__csr_mip__rg_usip$EN ; 
    reg RTL__csr_regfile__csr_mip__rg_utip ; 
    wire RTL__csr_regfile__csr_mip__rg_utip$D_IN , RTL__csr_regfile__csr_mip__rg_utip$EN ; 
    wire RTL__csr_regfile__csr_mip__CAN_FIRE_fav_write , RTL__csr_regfile__csr_mip__CAN_FIRE_m_external_interrupt_req , RTL__csr_regfile__csr_mip__CAN_FIRE_reset , RTL__csr_regfile__csr_mip__CAN_FIRE_s_external_interrupt_req , RTL__csr_regfile__csr_mip__CAN_FIRE_software_interrupt_req , RTL__csr_regfile__csr_mip__CAN_FIRE_timer_interrupt_req , RTL__csr_regfile__csr_mip__WILL_FIRE_fav_write , RTL__csr_regfile__csr_mip__WILL_FIRE_m_external_interrupt_req , RTL__csr_regfile__csr_mip__WILL_FIRE_reset , RTL__csr_regfile__csr_mip__WILL_FIRE_s_external_interrupt_req , RTL__csr_regfile__csr_mip__WILL_FIRE_software_interrupt_req , RTL__csr_regfile__csr_mip__WILL_FIRE_timer_interrupt_req ; 
    wire[11:0] RTL__csr_regfile__csr_mip__new_mip__h524 , RTL__csr_regfile__csr_mip__new_mip__h942 ; 
    wire RTL__csr_regfile__csr_mip__seip__h558 , RTL__csr_regfile__csr_mip__ssip__h562 , RTL__csr_regfile__csr_mip__stip__h560 , RTL__csr_regfile__csr_mip__ueip__h559 , RTL__csr_regfile__csr_mip__usip__h563 , RTL__csr_regfile__csr_mip__utip__h561 ; 
  assign  RTL__csr_regfile__csr_mip__CAN_FIRE_reset =1'd1; 
  assign  RTL__csr_regfile__csr_mip__WILL_FIRE_reset = RTL__csr_regfile__csr_mip__EN_reset ; 
  assign  RTL__csr_regfile__csr_mip__fv_read ={20'd0, RTL__csr_regfile__csr_mip__new_mip__h524 }; 
  assign  RTL__csr_regfile__csr_mip__fav_write ={20'd0, RTL__csr_regfile__csr_mip__new_mip__h942 }; 
  assign  RTL__csr_regfile__csr_mip__CAN_FIRE_fav_write =1'd1; 
  assign  RTL__csr_regfile__csr_mip__WILL_FIRE_fav_write = RTL__csr_regfile__csr_mip__EN_fav_write ; 
  assign  RTL__csr_regfile__csr_mip__CAN_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__WILL_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__CAN_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__WILL_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__CAN_FIRE_software_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__WILL_FIRE_software_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__CAN_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__WILL_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL__csr_regfile__csr_mip__rg_meip$D_IN = RTL__csr_regfile__csr_mip__m_external_interrupt_req_req ; 
  assign  RTL__csr_regfile__csr_mip__rg_meip$EN =1'b1; 
  assign  RTL__csr_regfile__csr_mip__rg_msip$D_IN = RTL__csr_regfile__csr_mip__software_interrupt_req_req ; 
  assign  RTL__csr_regfile__csr_mip__rg_msip$EN =1'b1; 
  assign  RTL__csr_regfile__csr_mip__rg_mtip$D_IN = RTL__csr_regfile__csr_mip__timer_interrupt_req_req ; 
  assign  RTL__csr_regfile__csr_mip__rg_mtip$EN =1'b1; 
  assign  RTL__csr_regfile__csr_mip__rg_seip$D_IN = RTL__csr_regfile__csr_mip__s_external_interrupt_req_req ; 
  assign  RTL__csr_regfile__csr_mip__rg_seip$EN =1'b1; 
  assign  RTL__csr_regfile__csr_mip__rg_ssip$D_IN =! RTL__csr_regfile__csr_mip__EN_reset && RTL__csr_regfile__csr_mip__ssip__h562 ; 
  assign  RTL__csr_regfile__csr_mip__rg_ssip$EN = RTL__csr_regfile__csr_mip__EN_fav_write || RTL__csr_regfile__csr_mip__EN_reset ; 
  assign  RTL__csr_regfile__csr_mip__rg_stip$D_IN =! RTL__csr_regfile__csr_mip__EN_reset && RTL__csr_regfile__csr_mip__stip__h560 ; 
  assign  RTL__csr_regfile__csr_mip__rg_stip$EN = RTL__csr_regfile__csr_mip__EN_fav_write || RTL__csr_regfile__csr_mip__EN_reset ; 
  assign  RTL__csr_regfile__csr_mip__rg_ueip$D_IN =! RTL__csr_regfile__csr_mip__EN_reset && RTL__csr_regfile__csr_mip__ueip__h559 ; 
  assign  RTL__csr_regfile__csr_mip__rg_ueip$EN = RTL__csr_regfile__csr_mip__EN_fav_write || RTL__csr_regfile__csr_mip__EN_reset ; 
  assign  RTL__csr_regfile__csr_mip__rg_usip$D_IN =! RTL__csr_regfile__csr_mip__EN_reset && RTL__csr_regfile__csr_mip__usip__h563 ; 
  assign  RTL__csr_regfile__csr_mip__rg_usip$EN = RTL__csr_regfile__csr_mip__EN_fav_write || RTL__csr_regfile__csr_mip__EN_reset ; 
  assign  RTL__csr_regfile__csr_mip__rg_utip$D_IN =! RTL__csr_regfile__csr_mip__EN_reset && RTL__csr_regfile__csr_mip__utip__h561 ; 
  assign  RTL__csr_regfile__csr_mip__rg_utip$EN = RTL__csr_regfile__csr_mip__EN_fav_write || RTL__csr_regfile__csr_mip__EN_reset ; 
  assign  RTL__csr_regfile__csr_mip__new_mip__h524 ={ RTL__csr_regfile__csr_mip__rg_meip ,1'b0, RTL__csr_regfile__csr_mip__rg_seip , RTL__csr_regfile__csr_mip__rg_ueip , RTL__csr_regfile__csr_mip__rg_mtip ,1'b0, RTL__csr_regfile__csr_mip__rg_stip , RTL__csr_regfile__csr_mip__rg_utip , RTL__csr_regfile__csr_mip__rg_msip ,1'b0, RTL__csr_regfile__csr_mip__rg_ssip , RTL__csr_regfile__csr_mip__rg_usip }; 
  assign  RTL__csr_regfile__csr_mip__new_mip__h942 ={ RTL__csr_regfile__csr_mip__rg_meip ,1'b0, RTL__csr_regfile__csr_mip__seip__h558 , RTL__csr_regfile__csr_mip__ueip__h559 , RTL__csr_regfile__csr_mip__rg_mtip ,1'b0, RTL__csr_regfile__csr_mip__stip__h560 , RTL__csr_regfile__csr_mip__utip__h561 , RTL__csr_regfile__csr_mip__rg_msip ,1'b0, RTL__csr_regfile__csr_mip__ssip__h562 , RTL__csr_regfile__csr_mip__usip__h563 }; 
  assign  RTL__csr_regfile__csr_mip__seip__h558 = RTL__csr_regfile__csr_mip__fav_write_misa [18]&& RTL__csr_regfile__csr_mip__fav_write_wordxl [9]; 
  assign  RTL__csr_regfile__csr_mip__ssip__h562 = RTL__csr_regfile__csr_mip__fav_write_misa [18]&& RTL__csr_regfile__csr_mip__fav_write_wordxl [1]; 
  assign  RTL__csr_regfile__csr_mip__stip__h560 = RTL__csr_regfile__csr_mip__fav_write_misa [18]&& RTL__csr_regfile__csr_mip__fav_write_wordxl [5]; 
  assign  RTL__csr_regfile__csr_mip__ueip__h559 = RTL__csr_regfile__csr_mip__fav_write_misa [13]&& RTL__csr_regfile__csr_mip__fav_write_wordxl [8]; 
  assign  RTL__csr_regfile__csr_mip__usip__h563 = RTL__csr_regfile__csr_mip__fav_write_misa [13]&& RTL__csr_regfile__csr_mip__fav_write_wordxl [0]; 
  assign  RTL__csr_regfile__csr_mip__utip__h561 = RTL__csr_regfile__csr_mip__fav_write_misa [13]&& RTL__csr_regfile__csr_mip__fav_write_wordxl [4]; 
  always @( posedge  RTL__csr_regfile__csr_mip__CLK )
         begin 
             if ( RTL__csr_regfile__csr_mip__RST_N ==1'b0)
                 begin  
                     RTL__csr_regfile__csr_mip__rg_meip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_msip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_mtip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_seip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_ssip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_stip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_ueip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_usip  <=1'd0; 
                     RTL__csr_regfile__csr_mip__rg_utip  <=1'd0;
                 end 
              else 
                 begin 
                     if ( RTL__csr_regfile__csr_mip__rg_meip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_meip  <= RTL__csr_regfile__csr_mip__rg_meip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_msip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_msip  <= RTL__csr_regfile__csr_mip__rg_msip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_mtip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_mtip  <= RTL__csr_regfile__csr_mip__rg_mtip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_seip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_seip  <= RTL__csr_regfile__csr_mip__rg_seip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_ssip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_ssip  <= RTL__csr_regfile__csr_mip__rg_ssip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_stip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_stip  <= RTL__csr_regfile__csr_mip__rg_stip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_ueip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_ueip  <= RTL__csr_regfile__csr_mip__rg_ueip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_usip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_usip  <= RTL__csr_regfile__csr_mip__rg_usip$D_IN ;
                     if ( RTL__csr_regfile__csr_mip__rg_utip$EN ) 
                         RTL__csr_regfile__csr_mip__rg_utip  <= RTL__csr_regfile__csr_mip__rg_utip$D_IN ;
                 end 
         end
 
    assign RTL__csr_regfile__csr_mip__CLK = RTL__csr_regfile__CLK;
    assign RTL__csr_regfile__csr_mip__RST_N = RTL__csr_regfile__RST_N;
    assign RTL__csr_regfile__csr_mip__EN_reset = RTL__csr_regfile__csr_mip$EN_reset;
    assign RTL__csr_regfile__csr_mip$fv_read = RTL__csr_regfile__csr_mip__fv_read;
    assign RTL__csr_regfile__csr_mip__fav_write_misa = RTL__csr_regfile__csr_mip$fav_write_misa;
    assign RTL__csr_regfile__csr_mip__fav_write_wordxl = RTL__csr_regfile__csr_mip$fav_write_wordxl;
    assign RTL__csr_regfile__csr_mip__EN_fav_write = RTL__csr_regfile__csr_mip$EN_fav_write;
    assign RTL__csr_regfile__csr_mip$fav_write = RTL__csr_regfile__csr_mip__fav_write;
    assign RTL__csr_regfile__csr_mip__m_external_interrupt_req_req = RTL__csr_regfile__csr_mip$m_external_interrupt_req_req;
    assign RTL__csr_regfile__csr_mip__s_external_interrupt_req_req = RTL__csr_regfile__csr_mip$s_external_interrupt_req_req;
    assign RTL__csr_regfile__csr_mip__software_interrupt_req_req = RTL__csr_regfile__csr_mip$software_interrupt_req_req;
    assign RTL__csr_regfile__csr_mip__timer_interrupt_req_req = RTL__csr_regfile__csr_mip$timer_interrupt_req_req;
      
    wire RTL__csr_regfile__f_reset_rsps__RST;
    wire RTL__csr_regfile__f_reset_rsps__CLK;
    wire RTL__csr_regfile__f_reset_rsps__ENQ;
    wire RTL__csr_regfile__f_reset_rsps__CLR;
    wire RTL__csr_regfile__f_reset_rsps__DEQ;
    wire RTL__csr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage1_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL__stage1_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL__stage1_f_reset_rsps__FULL_N;
    wire RTL__stage1_f_reset_rsps__EMPTY_N;
    wire RTL__stage1_f_reset_rsps__RST;
    wire RTL__stage1_f_reset_rsps__CLK;
    wire RTL__stage2_f_reset_reqs__ENQ;
    wire RTL__stage2_f_reset_reqs__CLR;
    wire RTL__stage2_f_reset_reqs__DEQ;
    wire RTL__stage2_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage2_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL__stage3_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL__stage3_f_reset_reqs__FULL_N;
    wire RTL__stage3_f_reset_reqs__EMPTY_N;
    wire RTL__stage3_f_reset_reqs__RST;
    wire RTL__stage3_f_reset_reqs__CLK;
    wire RTL__stage3_f_reset_reqs__ENQ;
    wire RTL__stage3_f_reset_reqs__CLR;
    wire RTL__stage3_f_reset_rsps__DEQ;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__stage3_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;

    parameter RTL__csr_regfile__f_reset_rsps__guarded =1; 
    reg RTL__csr_regfile__f_reset_rsps__empty_reg ; 
    reg RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__FULL_N = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__EMPTY_N = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__csr_regfile__f_reset_rsps__CLK )
         begin 
             if ( RTL__csr_regfile__f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__csr_regfile__f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__csr_regfile__f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__csr_regfile__f_reset_rsps__CLR )
                         begin  
                             RTL__csr_regfile__f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__csr_regfile__f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__csr_regfile__f_reset_rsps__ENQ &&! RTL__csr_regfile__f_reset_rsps__DEQ )
                             begin  
                                 RTL__csr_regfile__f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__csr_regfile__f_reset_rsps__full_reg  <=! RTL__csr_regfile__f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if (! RTL__csr_regfile__f_reset_rsps__ENQ && RTL__csr_regfile__f_reset_rsps__DEQ )
                                 begin  
                                     RTL__csr_regfile__f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__csr_regfile__f_reset_rsps__empty_reg  <=! RTL__csr_regfile__f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__csr_regfile__f_reset_rsps__CLK )
         begin : RTL__csr_regfile__f_reset_rsps__error_checks 
           reg RTL__csr_regfile__f_reset_rsps__deqerror , RTL__csr_regfile__f_reset_rsps__enqerror ; 
             RTL__csr_regfile__f_reset_rsps__deqerror  =0; 
             RTL__csr_regfile__f_reset_rsps__enqerror  =0;
             if ( RTL__csr_regfile__f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__csr_regfile__f_reset_rsps__empty_reg && RTL__csr_regfile__f_reset_rsps__DEQ )
                         begin  
                             RTL__csr_regfile__f_reset_rsps__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__csr_regfile__f_reset_rsps__full_reg && RTL__csr_regfile__f_reset_rsps__ENQ &&(! RTL__csr_regfile__f_reset_rsps__DEQ || RTL__csr_regfile__f_reset_rsps__guarded ))
                         begin  
                             RTL__csr_regfile__f_reset_rsps__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__csr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__empty_reg ;
      
    wire RTL__csr_regfile__soc_map__CLK;
    wire RTL__csr_regfile__soc_map__RST_N;
    wire[63:0] RTL__csr_regfile__soc_map__m_near_mem_io_addr_base;
    wire[63:0] RTL__csr_regfile__soc_map__m_near_mem_io_addr_size;
    wire[63:0] RTL__csr_regfile__soc_map__m_near_mem_io_addr_lim;
    wire[63:0] RTL__csr_regfile__soc_map__m_plic_addr_base;
    wire[63:0] RTL__csr_regfile__soc_map__m_plic_addr_size;
    wire[63:0] RTL__csr_regfile__soc_map__m_plic_addr_lim;
    wire[63:0] RTL__csr_regfile__soc_map__m_uart0_addr_base;
    wire[63:0] RTL__csr_regfile__soc_map__m_uart0_addr_size;
    wire[63:0] RTL__csr_regfile__soc_map__m_uart0_addr_lim;
    wire[63:0] RTL__csr_regfile__soc_map__m_boot_rom_addr_base;
    wire[63:0] RTL__csr_regfile__soc_map__m_boot_rom_addr_size;
    wire[63:0] RTL__csr_regfile__soc_map__m_boot_rom_addr_lim;
    wire[63:0] RTL__csr_regfile__soc_map__m_mem0_controller_addr_base;
    wire[63:0] RTL__csr_regfile__soc_map__m_mem0_controller_addr_size;
    wire[63:0] RTL__csr_regfile__soc_map__m_mem0_controller_addr_lim;
    wire[63:0] RTL__csr_regfile__soc_map__m_tcm_addr_base;
    wire[63:0] RTL__csr_regfile__soc_map__m_tcm_addr_size;
    wire[63:0] RTL__csr_regfile__soc_map__m_tcm_addr_lim;
    wire[63:0] RTL__csr_regfile__soc_map__m_is_mem_addr_addr;
    wire RTL__csr_regfile__soc_map__m_is_mem_addr;
    wire[63:0] RTL__csr_regfile__soc_map__m_is_IO_addr_addr;
    wire RTL__csr_regfile__soc_map__m_is_IO_addr;
    wire[63:0] RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr_addr;
    wire RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr;
    wire[63:0] RTL__csr_regfile__soc_map__m_pc_reset_value;
    wire[63:0] RTL__csr_regfile__soc_map__m_mtvec_reset_value;
    wire[63:0] RTL__csr_regfile__soc_map__m_nmivec_reset_value;
    wire RTL__soc_map__CLK;
    wire RTL__soc_map__RST_N;
    wire[63:0] RTL__soc_map__m_near_mem_io_addr_base;
    wire[63:0] RTL__soc_map__m_near_mem_io_addr_size;
    wire[63:0] RTL__soc_map__m_near_mem_io_addr_lim;
    wire[63:0] RTL__soc_map__m_plic_addr_base;
    wire[63:0] RTL__soc_map__m_plic_addr_size;
    wire[63:0] RTL__soc_map__m_plic_addr_lim;
    wire[63:0] RTL__soc_map__m_uart0_addr_base;
    wire[63:0] RTL__soc_map__m_uart0_addr_size;
    wire[63:0] RTL__soc_map__m_uart0_addr_lim;
    wire[63:0] RTL__soc_map__m_boot_rom_addr_base;
    wire[63:0] RTL__soc_map__m_boot_rom_addr_size;
    wire[63:0] RTL__soc_map__m_boot_rom_addr_lim;
    wire[63:0] RTL__soc_map__m_mem0_controller_addr_base;
    wire[63:0] RTL__soc_map__m_mem0_controller_addr_size;
    wire[63:0] RTL__soc_map__m_mem0_controller_addr_lim;
    wire[63:0] RTL__soc_map__m_tcm_addr_base;
    wire[63:0] RTL__soc_map__m_tcm_addr_size;
    wire[63:0] RTL__soc_map__m_tcm_addr_lim;
    wire[63:0] RTL__soc_map__m_is_mem_addr_addr;
    wire RTL__soc_map__m_is_mem_addr;
    wire[63:0] RTL__soc_map__m_is_IO_addr_addr;
    wire RTL__soc_map__m_is_IO_addr;
    wire[63:0] RTL__soc_map__m_is_near_mem_IO_addr_addr;
    wire RTL__soc_map__m_is_near_mem_IO_addr;
    wire[63:0] RTL__soc_map__m_pc_reset_value;
    wire[63:0] RTL__soc_map__m_mtvec_reset_value;
    wire[63:0] RTL__soc_map__m_nmivec_reset_value;

    wire[63:0] RTL__csr_regfile__soc_map__m_boot_rom_addr_base , RTL__csr_regfile__soc_map__m_boot_rom_addr_lim , RTL__csr_regfile__soc_map__m_boot_rom_addr_size , RTL__csr_regfile__soc_map__m_mem0_controller_addr_base , RTL__csr_regfile__soc_map__m_mem0_controller_addr_lim , RTL__csr_regfile__soc_map__m_mem0_controller_addr_size , RTL__csr_regfile__soc_map__m_mtvec_reset_value , RTL__csr_regfile__soc_map__m_near_mem_io_addr_base , RTL__csr_regfile__soc_map__m_near_mem_io_addr_lim , RTL__csr_regfile__soc_map__m_near_mem_io_addr_size , RTL__csr_regfile__soc_map__m_nmivec_reset_value , RTL__csr_regfile__soc_map__m_pc_reset_value , RTL__csr_regfile__soc_map__m_plic_addr_base , RTL__csr_regfile__soc_map__m_plic_addr_lim , RTL__csr_regfile__soc_map__m_plic_addr_size , RTL__csr_regfile__soc_map__m_tcm_addr_base , RTL__csr_regfile__soc_map__m_tcm_addr_lim , RTL__csr_regfile__soc_map__m_tcm_addr_size , RTL__csr_regfile__soc_map__m_uart0_addr_base , RTL__csr_regfile__soc_map__m_uart0_addr_lim , RTL__csr_regfile__soc_map__m_uart0_addr_size ; 
    wire RTL__csr_regfile__soc_map__m_is_IO_addr , RTL__csr_regfile__soc_map__m_is_mem_addr , RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr ; 
  assign  RTL__csr_regfile__soc_map__m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL__csr_regfile__soc_map__m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL__csr_regfile__soc_map__m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL__csr_regfile__soc_map__m_plic_addr_base =64'h000000000C000000; 
  assign  RTL__csr_regfile__soc_map__m_plic_addr_size =64'h0000000000400000; 
  assign  RTL__csr_regfile__soc_map__m_plic_addr_lim =64'd205520896; 
  assign  RTL__csr_regfile__soc_map__m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL__csr_regfile__soc_map__m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL__csr_regfile__soc_map__m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL__csr_regfile__soc_map__m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL__csr_regfile__soc_map__m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL__csr_regfile__soc_map__m_boot_rom_addr_lim =64'd8192; 
  assign  RTL__csr_regfile__soc_map__m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL__csr_regfile__soc_map__m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL__csr_regfile__soc_map__m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL__csr_regfile__soc_map__m_tcm_addr_base =64'h0; 
  assign  RTL__csr_regfile__soc_map__m_tcm_addr_size =64'd0; 
  assign  RTL__csr_regfile__soc_map__m_tcm_addr_lim =64'd0; 
  assign  RTL__csr_regfile__soc_map__m_is_mem_addr = RTL__csr_regfile__soc_map__m_is_mem_addr_addr >=64'h0000000000001000&& RTL__csr_regfile__soc_map__m_is_mem_addr_addr <64'd8192|| RTL__csr_regfile__soc_map__m_is_mem_addr_addr >=64'h0000000080000000&& RTL__csr_regfile__soc_map__m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL__csr_regfile__soc_map__m_is_IO_addr = RTL__csr_regfile__soc_map__m_is_IO_addr_addr >=64'h0000000002000000&& RTL__csr_regfile__soc_map__m_is_IO_addr_addr <64'd33603584|| RTL__csr_regfile__soc_map__m_is_IO_addr_addr >=64'h000000000C000000&& RTL__csr_regfile__soc_map__m_is_IO_addr_addr <64'd205520896|| RTL__csr_regfile__soc_map__m_is_IO_addr_addr >=64'h00000000C0000000&& RTL__csr_regfile__soc_map__m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr = RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL__csr_regfile__soc_map__m_pc_reset_value =64'h0000000000001000; 
  assign  RTL__csr_regfile__soc_map__m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL__csr_regfile__soc_map__m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
     
  assign  RTL__csr_regfile__CAN_FIRE_RL_rl_reset_start =! RTL__csr_regfile__rg_state ; 
  assign  RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start = RTL__csr_regfile__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__csr_regfile__CAN_FIRE_RL_rl_mcycle_incr =1'd1; 
  assign  RTL__csr_regfile__WILL_FIRE_RL_rl_mcycle_incr =1'd1; 
  assign  RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_csrrx = RTL__csr_regfile__MUX_rw_minstret$wset_1__SEL_1 || RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_csrrx = RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_csrrx ; 
  assign  RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_incr =! RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_csrrx && RTL__csr_regfile__EN_csr_minstret_incr ; 
  assign  RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_incr = RTL__csr_regfile__CAN_FIRE_RL_rl_upd_minstret_incr ; 
  assign  RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__SEL_2 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h300; 
  assign  RTL__csr_regfile__MUX_rg_mcause$write_1__SEL_2 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h342; 
  assign  RTL__csr_regfile__MUX_rg_mcounteren$write_1__SEL_1 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h306; 
  assign  RTL__csr_regfile__MUX_rg_mepc$write_1__SEL_1 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h341; 
  assign  RTL__csr_regfile__MUX_rg_mtval$write_1__SEL_1 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h343; 
  assign  RTL__csr_regfile__MUX_rg_mtvec$write_1__SEL_1 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h305; 
  assign  RTL__csr_regfile__MUX_rg_state$write_1__SEL_2 = RTL__csr_regfile__CAN_FIRE_RL_rl_reset_start &&! RTL__csr_regfile__EN_mav_csr_write ; 
  assign  RTL__csr_regfile__MUX_rg_tdata1$write_1__SEL_1 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h7A1; 
  assign  RTL__csr_regfile__MUX_rw_minstret$wset_1__SEL_1 = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d642 &&( RTL__csr_regfile__mav_csr_write_csr_addr ==12'hB02|| RTL__csr_regfile__mav_csr_write_csr_addr ==12'hB82); 
  assign  RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__VAL_3 ={9'd0, RTL__csr_regfile__fixed_up_val_23__h8130 }; 
  assign  RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_2 ={ RTL__csr_regfile__mav_csr_write_word [31], RTL__csr_regfile__mav_csr_write_word [3:0]}; 
  assign  RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_3 ={! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt , RTL__csr_regfile__exc_code__h7909 }; 
  assign  RTL__csr_regfile__MUX_rg_minstret$write_1__VAL_1 = RTL__csr_regfile__MUX_rw_minstret$wset_1__SEL_1  ?  RTL__csr_regfile__MUX_rw_minstret$wset_1__VAL_1 :64'd0; 
  assign  RTL__csr_regfile__MUX_rg_minstret$write_1__VAL_2 = RTL__csr_regfile__rg_minstret +64'd1; 
  assign  RTL__csr_regfile__MUX_rg_mtvec$write_1__VAL_1 ={ RTL__csr_regfile__mav_csr_write_word [31:2], RTL__csr_regfile__mav_csr_write_word [0]}; 
  assign  RTL__csr_regfile__MUX_rg_mtvec$write_1__VAL_2 ={ RTL__csr_regfile__soc_map$m_mtvec_reset_value [31:2], RTL__csr_regfile__soc_map$m_mtvec_reset_value [0]}; 
  assign  RTL__csr_regfile__MUX_rw_minstret$wset_1__VAL_1 =( RTL__csr_regfile__mav_csr_write_csr_addr ==12'hB02) ?  RTL__csr_regfile__x__h5174 : RTL__csr_regfile__x__h5282 ; 
  assign  RTL__csr_regfile__cfg_verbosity$D_IN =4'h0; 
  assign  RTL__csr_regfile__cfg_verbosity$EN =1'b0; 
  always @(        RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start                      or   RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__SEL_2               or   RTL__csr_regfile__wordxl1__h4038              or   RTL__csr_regfile__EN_csr_ret_actions             or   RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__VAL_3            or   RTL__csr_regfile__EN_csr_trap_actions           or   RTL__csr_regfile__x__h8067  )
         case (1'b1) 
          RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start  : 
              RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN  =32'd0; 
          RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__SEL_2  : 
              RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN  = RTL__csr_regfile__wordxl1__h4038 ; 
          RTL__csr_regfile__EN_csr_ret_actions  : 
              RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN  = RTL__csr_regfile__MUX_csr_mstatus_rg_mstatus$write_1__VAL_3 ; 
          RTL__csr_regfile__EN_csr_trap_actions  : 
              RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN  = RTL__csr_regfile__x__h8067 ;
          default : 
              RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN  =32'hAAAAAAAA;endcase
  assign  RTL__csr_regfile__csr_mstatus_rg_mstatus$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h300|| RTL__csr_regfile__EN_csr_trap_actions || RTL__csr_regfile__EN_csr_ret_actions || RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__rg_dcsr$D_IN =32'h0; 
  assign  RTL__csr_regfile__rg_dcsr$EN =1'b0; 
  assign  RTL__csr_regfile__rg_dpc$D_IN =32'h0; 
  assign  RTL__csr_regfile__rg_dpc$EN =1'b0; 
  assign  RTL__csr_regfile__rg_dscratch0$D_IN =32'h0; 
  assign  RTL__csr_regfile__rg_dscratch0$EN =1'b0; 
  assign  RTL__csr_regfile__rg_dscratch1$D_IN =32'h0; 
  assign  RTL__csr_regfile__rg_dscratch1$EN =1'b0; 
  always @(      RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start                  or   RTL__csr_regfile__MUX_rg_mcause$write_1__SEL_2             or   RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_2            or   RTL__csr_regfile__EN_csr_trap_actions           or   RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_3  )
         case (1'b1) 
          RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start  : 
              RTL__csr_regfile__rg_mcause$D_IN  =5'd0; 
          RTL__csr_regfile__MUX_rg_mcause$write_1__SEL_2  : 
              RTL__csr_regfile__rg_mcause$D_IN  = RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_2 ; 
          RTL__csr_regfile__EN_csr_trap_actions  : 
              RTL__csr_regfile__rg_mcause$D_IN  = RTL__csr_regfile__MUX_rg_mcause$write_1__VAL_3 ;
          default : 
              RTL__csr_regfile__rg_mcause$D_IN  =5'b01010;endcase
  assign  RTL__csr_regfile__rg_mcause$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h342|| RTL__csr_regfile__EN_csr_trap_actions || RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__rg_mcounteren$D_IN = RTL__csr_regfile__MUX_rg_mcounteren$write_1__SEL_1  ?  RTL__csr_regfile__mav_csr_write_word [2:0]:3'd0; 
  assign  RTL__csr_regfile__rg_mcounteren$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h306|| RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__rg_mcycle$D_IN = RTL__csr_regfile__rg_mcycle +64'd1; 
  assign  RTL__csr_regfile__rg_mcycle$EN =1'd1; 
  assign  RTL__csr_regfile__rg_mepc$D_IN = RTL__csr_regfile__MUX_rg_mepc$write_1__SEL_1  ?  RTL__csr_regfile__result__h4701 : RTL__csr_regfile__csr_trap_actions_pc ; 
  assign  RTL__csr_regfile__rg_mepc$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h341|| RTL__csr_regfile__EN_csr_trap_actions ; 
  assign  RTL__csr_regfile__rg_minstret$D_IN = RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_csrrx  ?  RTL__csr_regfile__MUX_rg_minstret$write_1__VAL_1 : RTL__csr_regfile__MUX_rg_minstret$write_1__VAL_2 ; 
  assign  RTL__csr_regfile__rg_minstret$EN = RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_csrrx || RTL__csr_regfile__WILL_FIRE_RL_rl_upd_minstret_incr ; 
  assign  RTL__csr_regfile__rg_mscratch$D_IN = RTL__csr_regfile__mav_csr_write_word ; 
  assign  RTL__csr_regfile__rg_mscratch$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h340; 
  assign  RTL__csr_regfile__rg_mtval$D_IN = RTL__csr_regfile__MUX_rg_mtval$write_1__SEL_1  ?  RTL__csr_regfile__mav_csr_write_word : RTL__csr_regfile__csr_trap_actions_xtval ; 
  assign  RTL__csr_regfile__rg_mtval$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h343|| RTL__csr_regfile__EN_csr_trap_actions ; 
  assign  RTL__csr_regfile__rg_mtvec$D_IN = RTL__csr_regfile__MUX_rg_mtvec$write_1__SEL_1  ?  RTL__csr_regfile__MUX_rg_mtvec$write_1__VAL_1 : RTL__csr_regfile__MUX_rg_mtvec$write_1__VAL_2 ; 
  assign  RTL__csr_regfile__rg_mtvec$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h305|| RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__rg_nmi$D_IN =! RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start && RTL__csr_regfile__nmi_req_set_not_clear ; 
  assign  RTL__csr_regfile__rg_nmi$EN =1'b1; 
  assign  RTL__csr_regfile__rg_nmi_vector$D_IN = RTL__csr_regfile__soc_map$m_nmivec_reset_value [31:0]; 
  assign  RTL__csr_regfile__rg_nmi_vector$EN = RTL__csr_regfile__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__csr_regfile__rg_state$D_IN =! RTL__csr_regfile__EN_server_reset_request_put ; 
  assign  RTL__csr_regfile__rg_state$EN = RTL__csr_regfile__EN_server_reset_request_put || RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__rg_tdata1$D_IN = RTL__csr_regfile__MUX_rg_tdata1$write_1__SEL_1  ?  RTL__csr_regfile__result__h5357 :32'd0; 
  assign  RTL__csr_regfile__rg_tdata1$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h7A1|| RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__rg_tdata2$D_IN = RTL__csr_regfile__mav_csr_write_word ; 
  assign  RTL__csr_regfile__rg_tdata2$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h7A2; 
  assign  RTL__csr_regfile__rg_tdata3$D_IN = RTL__csr_regfile__mav_csr_write_word ; 
  assign  RTL__csr_regfile__rg_tdata3$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h7A3; 
  assign  RTL__csr_regfile__rg_tselect$D_IN =32'd0; 
  assign  RTL__csr_regfile__rg_tselect$EN = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h7A0|| RTL__csr_regfile__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile__csr_mie$fav_write_misa =28'd68157696; 
  assign  RTL__csr_regfile__csr_mie$fav_write_wordxl = RTL__csr_regfile__mav_csr_write_word ; 
  assign  RTL__csr_regfile__csr_mie$EN_reset = RTL__csr_regfile__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__csr_regfile__csr_mie$EN_fav_write = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h304; 
  assign  RTL__csr_regfile__csr_mip$fav_write_misa =28'd68157696; 
  assign  RTL__csr_regfile__csr_mip$fav_write_wordxl = RTL__csr_regfile__mav_csr_write_word ; 
  assign  RTL__csr_regfile__csr_mip$m_external_interrupt_req_req = RTL__csr_regfile__m_external_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile__csr_mip$s_external_interrupt_req_req = RTL__csr_regfile__s_external_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile__csr_mip$software_interrupt_req_req = RTL__csr_regfile__software_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile__csr_mip$timer_interrupt_req_req = RTL__csr_regfile__timer_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile__csr_mip$EN_reset = RTL__csr_regfile__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__csr_regfile__csr_mip$EN_fav_write = RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL__csr_regfile__mav_csr_write_csr_addr ==12'h344; 
  assign  RTL__csr_regfile__f_reset_rsps$ENQ = RTL__csr_regfile__EN_server_reset_request_put ; 
  assign  RTL__csr_regfile__f_reset_rsps$DEQ = RTL__csr_regfile__EN_server_reset_response_get ; 
  assign  RTL__csr_regfile__f_reset_rsps$CLR =1'b0; 
  assign  RTL__csr_regfile__soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL__csr_regfile__soc_map$m_is_mem_addr_addr =64'h0; 
  assign  RTL__csr_regfile__soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1370 =(! RTL__csr_regfile__csr_mip$fv_read [11]||! RTL__csr_regfile__csr_mie$fv_read [11]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]) ? 4'd3:4'd11; 
  assign  RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1372 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339  ? 4'd9:( RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334  ? 4'd7: RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1370 ); 
  assign  RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1374 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349  ? 4'd5:( RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344  ? 4'd1: RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1372 ); 
  assign  RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1376 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359  ? 4'd0:( RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354  ? 4'd8: RTL__csr_regfile__IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1374 ); 
  assign  RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 =( RTL__csr_regfile__csr_ret_actions_from_priv ==2'b11) ?  RTL__csr_regfile___theResult___fst__h8211 : RTL__csr_regfile___theResult___fst__h8412 ; 
  assign  RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1068 =( RTL__csr_regfile__csr_ret_actions_from_priv ==2'b11) ? { RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [12:11], RTL__csr_regfile___theResult___fst__h8211 }:{ RTL__csr_regfile__to_y__h8411 , RTL__csr_regfile___theResult___fst__h8412 }; 
  assign  RTL__csr_regfile__NOT_access_permitted_1_csr_addr_ULT_0xC03_069__ETC___d1155 =( RTL__csr_regfile__access_permitted_1_csr_addr >=12'hC03&& RTL__csr_regfile__access_permitted_1_csr_addr <=12'hC1F|| RTL__csr_regfile__access_permitted_1_csr_addr >=12'hB03&& RTL__csr_regfile__access_permitted_1_csr_addr <=12'hB1F|| RTL__csr_regfile__access_permitted_1_csr_addr >=12'hC83&& RTL__csr_regfile__access_permitted_1_csr_addr <=12'hC9F|| RTL__csr_regfile__access_permitted_1_csr_addr >=12'hB83&& RTL__csr_regfile__access_permitted_1_csr_addr <=12'hB9F|| RTL__csr_regfile__access_permitted_1_csr_addr >=12'h323&& RTL__csr_regfile__access_permitted_1_csr_addr <=12'h33F|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hC00|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hC02|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hC80|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hC81|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hC82|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hF11|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hF12|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hF13|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hF14|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h300|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h301|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h304|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h305|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h306|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h340|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h341|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h342|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h343|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h344|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hB00|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hB02|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hB80|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'hB82|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h7A0|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h7A1|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h7A2|| RTL__csr_regfile__access_permitted_1_csr_addr ==12'h7A3)&& RTL__csr_regfile__access_permitted_1_priv >= RTL__csr_regfile__access_permitted_1_csr_addr [9:8]&&( RTL__csr_regfile__access_permitted_1_csr_addr !=12'h180||! RTL__csr_regfile__csr_mstatus_rg_mstatus [20]); 
  assign  RTL__csr_regfile__NOT_access_permitted_2_csr_addr_ULT_0xC03_160__ETC___d1245 =( RTL__csr_regfile__access_permitted_2_csr_addr >=12'hC03&& RTL__csr_regfile__access_permitted_2_csr_addr <=12'hC1F|| RTL__csr_regfile__access_permitted_2_csr_addr >=12'hB03&& RTL__csr_regfile__access_permitted_2_csr_addr <=12'hB1F|| RTL__csr_regfile__access_permitted_2_csr_addr >=12'hC83&& RTL__csr_regfile__access_permitted_2_csr_addr <=12'hC9F|| RTL__csr_regfile__access_permitted_2_csr_addr >=12'hB83&& RTL__csr_regfile__access_permitted_2_csr_addr <=12'hB9F|| RTL__csr_regfile__access_permitted_2_csr_addr >=12'h323&& RTL__csr_regfile__access_permitted_2_csr_addr <=12'h33F|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hC00|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hC02|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hC80|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hC81|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hC82|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hF11|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hF12|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hF13|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hF14|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h300|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h301|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h304|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h305|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h306|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h340|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h341|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h342|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h343|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h344|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hB00|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hB02|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hB80|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'hB82|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h7A0|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h7A1|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h7A2|| RTL__csr_regfile__access_permitted_2_csr_addr ==12'h7A3)&& RTL__csr_regfile__access_permitted_2_priv >= RTL__csr_regfile__access_permitted_2_csr_addr [9:8]&&( RTL__csr_regfile__access_permitted_2_csr_addr !=12'h180||! RTL__csr_regfile__csr_mstatus_rg_mstatus [20]); 
  assign  RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 = RTL__csr_regfile__cfg_verbosity >4'd1; 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334 =(! RTL__csr_regfile__csr_mip$fv_read [11]||! RTL__csr_regfile__csr_mie$fv_read [11]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3])&&(! RTL__csr_regfile__csr_mip$fv_read [3]||! RTL__csr_regfile__csr_mie$fv_read [3]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334 &&(! RTL__csr_regfile__csr_mip$fv_read [7]||! RTL__csr_regfile__csr_mie$fv_read [7]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339 &&(! RTL__csr_regfile__csr_mip$fv_read [9]||! RTL__csr_regfile__csr_mie$fv_read [9]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344 &&(! RTL__csr_regfile__csr_mip$fv_read [1]||! RTL__csr_regfile__csr_mie$fv_read [1]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349 &&(! RTL__csr_regfile__csr_mip$fv_read [5]||! RTL__csr_regfile__csr_mie$fv_read [5]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354 &&(! RTL__csr_regfile__csr_mip$fv_read [8]||! RTL__csr_regfile__csr_mie$fv_read [8]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1364 = RTL__csr_regfile__NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359 &&(! RTL__csr_regfile__csr_mip$fv_read [0]||! RTL__csr_regfile__csr_mie$fv_read [0]|| RTL__csr_regfile__interrupt_pending_cur_priv ==2'b11&&! RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__NOT_csr_trap_actions_nmi_97_AND_csr_trap_actio_ETC___d974 =! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 !=4'd0&& RTL__csr_regfile__exc_code__h7909 !=4'd1&& RTL__csr_regfile__exc_code__h7909 !=4'd2&& RTL__csr_regfile__exc_code__h7909 !=4'd3&& RTL__csr_regfile__exc_code__h7909 !=4'd4&& RTL__csr_regfile__exc_code__h7909 !=4'd5&& RTL__csr_regfile__exc_code__h7909 !=4'd6&& RTL__csr_regfile__exc_code__h7909 !=4'd7&& RTL__csr_regfile__exc_code__h7909 !=4'd8&& RTL__csr_regfile__exc_code__h7909 !=4'd9&& RTL__csr_regfile__exc_code__h7909 !=4'd10&& RTL__csr_regfile__exc_code__h7909 !=4'd11; 
  assign  RTL__csr_regfile__NOT_mav_csr_write_csr_addr_ULT_0xB03_77_35_AND_ETC___d746 =! RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03___d577 && RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB1F___d578 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB83___d581 && RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB9F___d582 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323___d585 && RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0x33F___d586 || RTL__csr_regfile__mav_csr_write_csr_addr ==12'hF11|| RTL__csr_regfile__mav_csr_write_csr_addr ==12'hF12|| RTL__csr_regfile__mav_csr_write_csr_addr ==12'hF13|| RTL__csr_regfile__mav_csr_write_csr_addr ==12'hF14; 
  assign  RTL__csr_regfile___theResult___fst__h8211 ={ RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [31:13],2'd0, RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [10:0]}; 
  assign  RTL__csr_regfile___theResult___fst__h8412 ={ RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [31:9],1'd0, RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [7:0]}; 
  assign  RTL__csr_regfile__b__h8248 = RTL__csr_regfile__csr_mstatus_rg_mstatus [{3'd1, RTL__csr_regfile__csr_ret_actions_from_priv }]; 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1288 = RTL__csr_regfile__csr_mip$fv_read [11]&& RTL__csr_regfile__csr_mie$fv_read [11]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3])|| RTL__csr_regfile__csr_mip$fv_read [3]&& RTL__csr_regfile__csr_mie$fv_read [3]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1293 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1288 || RTL__csr_regfile__csr_mip$fv_read [7]&& RTL__csr_regfile__csr_mie$fv_read [7]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1298 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1293 || RTL__csr_regfile__csr_mip$fv_read [9]&& RTL__csr_regfile__csr_mie$fv_read [9]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1303 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1298 || RTL__csr_regfile__csr_mip$fv_read [1]&& RTL__csr_regfile__csr_mie$fv_read [1]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1308 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1303 || RTL__csr_regfile__csr_mip$fv_read [5]&& RTL__csr_regfile__csr_mie$fv_read [5]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1313 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1308 || RTL__csr_regfile__csr_mip$fv_read [8]&& RTL__csr_regfile__csr_mie$fv_read [8]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1318 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1313 || RTL__csr_regfile__csr_mip$fv_read [0]&& RTL__csr_regfile__csr_mie$fv_read [0]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1323 = RTL__csr_regfile__csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1318 || RTL__csr_regfile__csr_mip$fv_read [4]&& RTL__csr_regfile__csr_mie$fv_read [4]&&( RTL__csr_regfile__interrupt_pending_cur_priv !=2'b11|| RTL__csr_regfile__csr_mstatus_rg_mstatus [3]); 
  assign  RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 = RTL__csr_regfile__x__h8244 | RTL__csr_regfile__mask__h8232 ; 
  assign  RTL__csr_regfile__csr_trap_actions_nmi_OR_NOT_csr_trap_actions_i_ETC___d1025 =( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 !=4'd0&& RTL__csr_regfile__exc_code__h7909 !=4'd1&& RTL__csr_regfile__exc_code__h7909 !=4'd2&& RTL__csr_regfile__exc_code__h7909 !=4'd3&& RTL__csr_regfile__exc_code__h7909 !=4'd4&& RTL__csr_regfile__exc_code__h7909 !=4'd5&& RTL__csr_regfile__exc_code__h7909 !=4'd6&& RTL__csr_regfile__exc_code__h7909 !=4'd7&& RTL__csr_regfile__exc_code__h7909 !=4'd8&& RTL__csr_regfile__exc_code__h7909 !=4'd9&& RTL__csr_regfile__exc_code__h7909 !=4'd11&& RTL__csr_regfile__exc_code__h7909 !=4'd12&& RTL__csr_regfile__exc_code__h7909 !=4'd13&& RTL__csr_regfile__exc_code__h7909 !=4'd15; 
  assign  RTL__csr_regfile__exc_code__h7909 = RTL__csr_regfile__csr_trap_actions_nmi  ? 4'd0: RTL__csr_regfile__csr_trap_actions_exc_code ; 
  assign  RTL__csr_regfile__exc_pc___1__h7296 = RTL__csr_regfile__exc_pc__h7243 + RTL__csr_regfile__vector_offset__h7244 ; 
  assign  RTL__csr_regfile__exc_pc__h7032 ={ RTL__csr_regfile__rg_mtvec [30:1],2'd0}; 
  assign  RTL__csr_regfile__exc_pc__h7243 = RTL__csr_regfile__csr_trap_actions_nmi  ?  RTL__csr_regfile__rg_nmi_vector : RTL__csr_regfile__exc_pc__h7032 ; 
  assign  RTL__csr_regfile__fixed_up_val_23__h4079 ={ RTL__csr_regfile__mav_csr_write_word [22:17],4'd0,( RTL__csr_regfile__mav_csr_write_word [12:11]==2'b11) ?  RTL__csr_regfile__mav_csr_write_word [12:11]:2'b0, RTL__csr_regfile__mav_csr_write_word [10:9],1'd0, RTL__csr_regfile__mav_csr_write_word [7:6],2'd0, RTL__csr_regfile__mav_csr_write_word [3:2],2'd0}; 
  assign  RTL__csr_regfile__fixed_up_val_23__h6471 ={ RTL__csr_regfile__csr_mstatus_rg_mstatus [22:17],4'd0, RTL__csr_regfile__mpp__h7337 , RTL__csr_regfile__csr_mstatus_rg_mstatus [10:9],1'd0, RTL__csr_regfile__csr_mstatus_rg_mstatus [3], RTL__csr_regfile__csr_mstatus_rg_mstatus [6],3'd0, RTL__csr_regfile__csr_mstatus_rg_mstatus [2],2'd0}; 
  assign  RTL__csr_regfile__fixed_up_val_23__h8130 ={ RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [22:17],4'd0,( RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [12:11]==2'b11) ?  RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [12:11]:2'b0, RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [10:9],1'd0, RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [7:6],2'd0, RTL__csr_regfile__IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [3:2],2'd0}; 
  assign  RTL__csr_regfile__ie_from_x__h8195 ={4'd0, RTL__csr_regfile__csr_ret_actions_from_priv }; 
  assign  RTL__csr_regfile__mask__h8232 =32'd1<< RTL__csr_regfile__pie_from_x__h8196 ; 
  assign  RTL__csr_regfile__mask__h8249 =32'd1<< RTL__csr_regfile__ie_from_x__h8195 ; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0x33F___d586 = RTL__csr_regfile__mav_csr_write_csr_addr <=12'h33F; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB1F___d578 = RTL__csr_regfile__mav_csr_write_csr_addr <=12'hB1F; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB9F___d582 = RTL__csr_regfile__mav_csr_write_csr_addr <=12'hB9F; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323_85_OR_NOT_mav_ETC___d728 =( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323___d585 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0x33F___d586 )&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF11&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF12&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF13&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF14&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h300&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h301&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h304&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h305&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h306&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h340&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h341&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h342&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h343&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h344&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hB00&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hB02&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hB80&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hB82&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h7A0&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h7A1&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h7A2&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'h7A3; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323___d585 = RTL__csr_regfile__mav_csr_write_csr_addr <12'h323; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 =( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03___d577 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB1F___d578 )&&( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB83___d581 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB9F___d582 )&&( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323___d585 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0x33F___d586 ); 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d642 =( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03___d577 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB1F___d578 )&&( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB83___d581 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB9F___d582 )&&( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323___d585 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0x33F___d586 )&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF11&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF12&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF13&& RTL__csr_regfile__mav_csr_write_csr_addr !=12'hF14; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d730 =( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03___d577 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB1F___d578 )&&( RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB83___d581 ||! RTL__csr_regfile__mav_csr_write_csr_addr_ULE_0xB9F___d582 )&& RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0x323_85_OR_NOT_mav_ETC___d728 ; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03___d577 = RTL__csr_regfile__mav_csr_write_csr_addr <12'hB03; 
  assign  RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB83___d581 = RTL__csr_regfile__mav_csr_write_csr_addr <12'hB83; 
  assign  RTL__csr_regfile__mpp__h7337 =( RTL__csr_regfile__csr_trap_actions_from_priv ==2'b11) ?  RTL__csr_regfile__csr_trap_actions_from_priv :2'b0; 
  assign  RTL__csr_regfile__pie_from_x__h8196 ={4'd1, RTL__csr_regfile__csr_ret_actions_from_priv }; 
  assign  RTL__csr_regfile__result__h4701 ={ RTL__csr_regfile__mav_csr_write_word [31:2],2'd0}; 
  assign  RTL__csr_regfile__result__h5357 ={4'd0, RTL__csr_regfile__mav_csr_write_word [27:0]}; 
  assign  RTL__csr_regfile__to_y__h8411 ={1'b0, RTL__csr_regfile__csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [8]}; 
  assign  RTL__csr_regfile__v__h4509 ={ RTL__csr_regfile__mav_csr_write_word [31:2],1'b0, RTL__csr_regfile__mav_csr_write_word [0]}; 
  assign  RTL__csr_regfile__v__h4571 ={29'd0, RTL__csr_regfile__mav_csr_write_word [2:0]}; 
  assign  RTL__csr_regfile__v__h4742 ={ RTL__csr_regfile__mav_csr_write_word [31],27'd0, RTL__csr_regfile__mav_csr_write_word [3:0]}; 
  assign  RTL__csr_regfile__val__h8250 ={31'd0, RTL__csr_regfile__b__h8248 }<< RTL__csr_regfile__ie_from_x__h8195 ; 
  assign  RTL__csr_regfile__vector_offset__h7244 ={26'd0, RTL__csr_regfile__csr_trap_actions_exc_code ,2'd0}; 
  assign  RTL__csr_regfile__wordxl1__h4038 ={9'd0, RTL__csr_regfile__fixed_up_val_23__h4079 }; 
  assign  RTL__csr_regfile__x__h5174 ={ RTL__csr_regfile__rg_minstret [63:32], RTL__csr_regfile__mav_csr_write_word }; 
  assign  RTL__csr_regfile__x__h5282 ={ RTL__csr_regfile__mav_csr_write_word , RTL__csr_regfile__rg_minstret [31:0]}; 
  assign  RTL__csr_regfile__x__h5843 =( RTL__csr_regfile__csr_trap_actions_interrupt &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__rg_mtvec [0]) ?  RTL__csr_regfile__exc_pc___1__h7296 : RTL__csr_regfile__exc_pc__h7243 ; 
  assign  RTL__csr_regfile__x__h8067 ={9'd0, RTL__csr_regfile__fixed_up_val_23__h6471 }; 
  assign  RTL__csr_regfile__x__h8068 ={! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt ,27'd0, RTL__csr_regfile__exc_code__h7909 }; 
  assign  RTL__csr_regfile__x__h8085 ={ RTL__csr_regfile__rg_mepc [31:2],1'd0, RTL__csr_regfile__rg_mepc [0]}; 
  assign  RTL__csr_regfile__x__h8231 = RTL__csr_regfile__x__h8261 | RTL__csr_regfile__val__h8250 ; 
  assign  RTL__csr_regfile__x__h8244 = RTL__csr_regfile__x__h8231 & RTL__csr_regfile__y__h8245 ; 
  assign  RTL__csr_regfile__x__h8261 = RTL__csr_regfile__csr_mstatus_rg_mstatus & RTL__csr_regfile__y__h8262 ; 
  assign  RTL__csr_regfile__y__h8245 =~ RTL__csr_regfile__mask__h8232 ; 
  assign  RTL__csr_regfile__y__h8262 =~ RTL__csr_regfile__mask__h8249 ; 
  always @(                 RTL__csr_regfile__read_csr_csr_addr                                        or   RTL__csr_regfile__rg_tdata3                        or   RTL__csr_regfile__csr_mstatus_rg_mstatus                       or   RTL__csr_regfile__csr_mie$fv_read                      or   RTL__csr_regfile__rg_mtvec                     or   RTL__csr_regfile__rg_mcounteren                    or   RTL__csr_regfile__rg_mscratch                   or   RTL__csr_regfile__x__h8085                  or   RTL__csr_regfile__rg_mcause                 or   RTL__csr_regfile__rg_mtval                or   RTL__csr_regfile__csr_mip$fv_read               or   RTL__csr_regfile__rg_tselect              or   RTL__csr_regfile__rg_tdata1             or   RTL__csr_regfile__rg_tdata2            or   RTL__csr_regfile__rg_mcycle           or   RTL__csr_regfile__rg_minstret  )
         begin 
             case ( RTL__csr_regfile__read_csr_csr_addr )
              12 'h300: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__csr_mstatus_rg_mstatus ;
              12 'h301: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  =32'd1074790656;
              12 'h304: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__csr_mie$fv_read ;
              12 'h305: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  ={ RTL__csr_regfile__rg_mtvec [30:1],1'b0, RTL__csr_regfile__rg_mtvec [0]};
              12 'h306: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  ={29'd0, RTL__csr_regfile__rg_mcounteren };
              12 'h340: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_mscratch ;
              12 'h341: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__x__h8085 ;
              12 'h342: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  ={ RTL__csr_regfile__rg_mcause [4],27'd0, RTL__csr_regfile__rg_mcause [3:0]};
              12 'h343: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_mtval ;
              12 'h344: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__csr_mip$fv_read ;
              12 'h7A0: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_tselect ;
              12 'h7A1: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_tdata1 ;
              12 'h7A2: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_tdata2 ;
              12 'hB00,12'hC00: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_mcycle [31:0];
              12 'hB02,12'hC02: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_minstret [31:0];
              12 'hB80,12'hC80: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_mcycle [63:32];
              12 'hB82,12'hC82: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_minstret [63:32];
              12 'hF11,12'hF12,12'hF13,12'hF14: 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  =32'd0;
              default : 
                  RTL__csr_regfile__IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL__csr_regfile__rg_tdata3 ;endcase
         end
  always @(                 RTL__csr_regfile__read_csr_port2_csr_addr                                        or   RTL__csr_regfile__rg_tdata3                        or   RTL__csr_regfile__csr_mstatus_rg_mstatus                       or   RTL__csr_regfile__csr_mie$fv_read                      or   RTL__csr_regfile__rg_mtvec                     or   RTL__csr_regfile__rg_mcounteren                    or   RTL__csr_regfile__rg_mscratch                   or   RTL__csr_regfile__x__h8085                  or   RTL__csr_regfile__rg_mcause                 or   RTL__csr_regfile__rg_mtval                or   RTL__csr_regfile__csr_mip$fv_read               or   RTL__csr_regfile__rg_tselect              or   RTL__csr_regfile__rg_tdata1             or   RTL__csr_regfile__rg_tdata2            or   RTL__csr_regfile__rg_mcycle           or   RTL__csr_regfile__rg_minstret  )
         begin 
             case ( RTL__csr_regfile__read_csr_port2_csr_addr )
              12 'h300: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__csr_mstatus_rg_mstatus ;
              12 'h301: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  =32'd1074790656;
              12 'h304: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__csr_mie$fv_read ;
              12 'h305: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  ={ RTL__csr_regfile__rg_mtvec [30:1],1'b0, RTL__csr_regfile__rg_mtvec [0]};
              12 'h306: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  ={29'd0, RTL__csr_regfile__rg_mcounteren };
              12 'h340: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_mscratch ;
              12 'h341: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__x__h8085 ;
              12 'h342: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  ={ RTL__csr_regfile__rg_mcause [4],27'd0, RTL__csr_regfile__rg_mcause [3:0]};
              12 'h343: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_mtval ;
              12 'h344: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__csr_mip$fv_read ;
              12 'h7A0: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_tselect ;
              12 'h7A1: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_tdata1 ;
              12 'h7A2: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_tdata2 ;
              12 'hB00,12'hC00: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_mcycle [31:0];
              12 'hB02,12'hC02: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_minstret [31:0];
              12 'hB80,12'hC80: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_mcycle [63:32];
              12 'hB82,12'hC82: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_minstret [63:32];
              12 'hF11,12'hF12,12'hF13,12'hF14: 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  =32'd0;
              default : 
                  RTL__csr_regfile__IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL__csr_regfile__rg_tdata3 ;endcase
         end
  always @(                 RTL__csr_regfile__mav_read_csr_csr_addr                                        or   RTL__csr_regfile__rg_tdata3                        or   RTL__csr_regfile__csr_mstatus_rg_mstatus                       or   RTL__csr_regfile__csr_mie$fv_read                      or   RTL__csr_regfile__rg_mtvec                     or   RTL__csr_regfile__rg_mcounteren                    or   RTL__csr_regfile__rg_mscratch                   or   RTL__csr_regfile__x__h8085                  or   RTL__csr_regfile__rg_mcause                 or   RTL__csr_regfile__rg_mtval                or   RTL__csr_regfile__csr_mip$fv_read               or   RTL__csr_regfile__rg_tselect              or   RTL__csr_regfile__rg_tdata1             or   RTL__csr_regfile__rg_tdata2            or   RTL__csr_regfile__rg_mcycle           or   RTL__csr_regfile__rg_minstret  )
         begin 
             case ( RTL__csr_regfile__mav_read_csr_csr_addr )
              12 'h300: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__csr_mstatus_rg_mstatus ;
              12 'h301: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  =32'd1074790656;
              12 'h304: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__csr_mie$fv_read ;
              12 'h305: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  ={ RTL__csr_regfile__rg_mtvec [30:1],1'b0, RTL__csr_regfile__rg_mtvec [0]};
              12 'h306: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  ={29'd0, RTL__csr_regfile__rg_mcounteren };
              12 'h340: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_mscratch ;
              12 'h341: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__x__h8085 ;
              12 'h342: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  ={ RTL__csr_regfile__rg_mcause [4],27'd0, RTL__csr_regfile__rg_mcause [3:0]};
              12 'h343: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_mtval ;
              12 'h344: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__csr_mip$fv_read ;
              12 'h7A0: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_tselect ;
              12 'h7A1: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_tdata1 ;
              12 'h7A2: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_tdata2 ;
              12 'hB00,12'hC00: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_mcycle [31:0];
              12 'hB02,12'hC02: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_minstret [31:0];
              12 'hB80,12'hC80: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_mcycle [63:32];
              12 'hB82,12'hC82: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_minstret [63:32];
              12 'hF11,12'hF12,12'hF13,12'hF14: 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  =32'd0;
              default : 
                  RTL__csr_regfile__IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL__csr_regfile__rg_tdata3 ;endcase
         end
  always @(           RTL__csr_regfile__mav_csr_write_csr_addr                            or   RTL__csr_regfile__mav_csr_write_word                  or   RTL__csr_regfile__wordxl1__h4038                 or   RTL__csr_regfile__csr_mie$fav_write                or   RTL__csr_regfile__v__h4509               or   RTL__csr_regfile__v__h4571              or   RTL__csr_regfile__result__h4701             or   RTL__csr_regfile__v__h4742            or   RTL__csr_regfile__csr_mip$fav_write           or   RTL__csr_regfile__result__h5357  )
         begin 
             case ( RTL__csr_regfile__mav_csr_write_csr_addr )
              12 'h300: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__wordxl1__h4038 ;
              12 'h301: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  =32'd1074790656;
              12 'h304: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__csr_mie$fav_write ;
              12 'h305: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__v__h4509 ;
              12 'h306: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__v__h4571 ;
              12 'h340,12'h343,12'hB00,12'hB02,12'hB80,12'hB82: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__mav_csr_write_word ;
              12 'h341: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__result__h4701 ;
              12 'h342: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__v__h4742 ;
              12 'h344: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__csr_mip$fav_write ;
              12 'h7A0: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  =32'd0;
              12 'h7A1: 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__result__h5357 ;
              default : 
                  RTL__csr_regfile__IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL__csr_regfile__mav_csr_write_word ;endcase
         end
  always @( posedge  RTL__csr_regfile__CLK )
         begin 
             if ( RTL__csr_regfile__RST_N ==1'b0)
                 begin  
                     RTL__csr_regfile__cfg_verbosity  <=4'd0; 
                     RTL__csr_regfile__csr_mstatus_rg_mstatus  <=32'd0; 
                     RTL__csr_regfile__rg_mcycle  <=64'd0; 
                     RTL__csr_regfile__rg_minstret  <=64'd0; 
                     RTL__csr_regfile__rg_nmi  <=1'd0; 
                     RTL__csr_regfile__rg_state  <=1'd0;
                 end 
              else 
                 begin 
                     if ( RTL__csr_regfile__cfg_verbosity$EN ) 
                         RTL__csr_regfile__cfg_verbosity  <= RTL__csr_regfile__cfg_verbosity$D_IN ;
                     if ( RTL__csr_regfile__csr_mstatus_rg_mstatus$EN ) 
                         RTL__csr_regfile__csr_mstatus_rg_mstatus  <= RTL__csr_regfile__csr_mstatus_rg_mstatus$D_IN ;
                     if ( RTL__csr_regfile__rg_mcycle$EN ) 
                         RTL__csr_regfile__rg_mcycle  <= RTL__csr_regfile__rg_mcycle$D_IN ;
                     if ( RTL__csr_regfile__rg_minstret$EN ) 
                         RTL__csr_regfile__rg_minstret  <= RTL__csr_regfile__rg_minstret$D_IN ;
                     if ( RTL__csr_regfile__rg_nmi$EN ) 
                         RTL__csr_regfile__rg_nmi  <= RTL__csr_regfile__rg_nmi$D_IN ;
                     if ( RTL__csr_regfile__rg_state$EN ) 
                         RTL__csr_regfile__rg_state  <= RTL__csr_regfile__rg_state$D_IN ;
                 end 
             if ( RTL__csr_regfile__rg_dcsr$EN ) 
                 RTL__csr_regfile__rg_dcsr  <= RTL__csr_regfile__rg_dcsr$D_IN ;
             if ( RTL__csr_regfile__rg_dpc$EN ) 
                 RTL__csr_regfile__rg_dpc  <= RTL__csr_regfile__rg_dpc$D_IN ;
             if ( RTL__csr_regfile__rg_dscratch0$EN ) 
                 RTL__csr_regfile__rg_dscratch0  <= RTL__csr_regfile__rg_dscratch0$D_IN ;
             if ( RTL__csr_regfile__rg_dscratch1$EN ) 
                 RTL__csr_regfile__rg_dscratch1  <= RTL__csr_regfile__rg_dscratch1$D_IN ;
             if ( RTL__csr_regfile__rg_mcause$EN ) 
                 RTL__csr_regfile__rg_mcause  <= RTL__csr_regfile__rg_mcause$D_IN ;
             if ( RTL__csr_regfile__rg_mcounteren$EN ) 
                 RTL__csr_regfile__rg_mcounteren  <= RTL__csr_regfile__rg_mcounteren$D_IN ;
             if ( RTL__csr_regfile__rg_mepc$EN ) 
                 RTL__csr_regfile__rg_mepc  <= RTL__csr_regfile__rg_mepc$D_IN ;
             if ( RTL__csr_regfile__rg_mscratch$EN ) 
                 RTL__csr_regfile__rg_mscratch  <= RTL__csr_regfile__rg_mscratch$D_IN ;
             if ( RTL__csr_regfile__rg_mtval$EN ) 
                 RTL__csr_regfile__rg_mtval  <= RTL__csr_regfile__rg_mtval$D_IN ;
             if ( RTL__csr_regfile__rg_mtvec$EN ) 
                 RTL__csr_regfile__rg_mtvec  <= RTL__csr_regfile__rg_mtvec$D_IN ;
             if ( RTL__csr_regfile__rg_nmi_vector$EN ) 
                 RTL__csr_regfile__rg_nmi_vector  <= RTL__csr_regfile__rg_nmi_vector$D_IN ;
             if ( RTL__csr_regfile__rg_tdata1$EN ) 
                 RTL__csr_regfile__rg_tdata1  <= RTL__csr_regfile__rg_tdata1$D_IN ;
             if ( RTL__csr_regfile__rg_tdata2$EN ) 
                 RTL__csr_regfile__rg_tdata2  <= RTL__csr_regfile__rg_tdata2$D_IN ;
             if ( RTL__csr_regfile__rg_tdata3$EN ) 
                 RTL__csr_regfile__rg_tdata3  <= RTL__csr_regfile__rg_tdata3$D_IN ;
             if ( RTL__csr_regfile__rg_tselect$EN ) 
                 RTL__csr_regfile__rg_tselect  <= RTL__csr_regfile__rg_tselect$D_IN ;
         end
  always @( negedge  RTL__csr_regfile__CLK )
         begin #0;
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_debug )$display("mstatus = 0x%0h", RTL__csr_regfile__csr_mstatus_rg_mstatus );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_debug )$display("mip     = 0x%0h", RTL__csr_regfile__csr_mip$fv_read );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_debug )$display("mie     = 0x%0h", RTL__csr_regfile__csr_mie$fv_read );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_Regfile.csr_trap_actions:", RTL__csr_regfile__rg_mcycle );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("    from priv %0d  pc 0x%0h  interrupt %0d  exc_code %0d  xtval 0x%0h", RTL__csr_regfile__csr_trap_actions_from_priv , RTL__csr_regfile__csr_trap_actions_pc , RTL__csr_regfile__csr_trap_actions_interrupt , RTL__csr_regfile__csr_trap_actions_exc_code , RTL__csr_regfile__csr_trap_actions_xtval );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("    priv %0d: ",2'b11);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ip: 0x%0h", RTL__csr_regfile__csr_mip$fv_read );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ie: 0x%0h", RTL__csr_regfile__csr_mie$fv_read );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" edeleg: 0x%0h",16'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ideleg: 0x%0h",12'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" cause:");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd0)$write("USER_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd1)$write("SUPERVISOR_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd2)$write("HYPERVISOR_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd3)$write("MACHINE_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd4)$write("USER_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd5)$write("SUPERVISOR_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd6)$write("HYPERVISOR_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd7)$write("MACHINE_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd8)$write("USER_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd9)$write("SUPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd10)$write("HYPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd11)$write("MACHINE_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]!=4'd0&& RTL__csr_regfile__rg_mcause [3:0]!=4'd1&& RTL__csr_regfile__rg_mcause [3:0]!=4'd2&& RTL__csr_regfile__rg_mcause [3:0]!=4'd3&& RTL__csr_regfile__rg_mcause [3:0]!=4'd4&& RTL__csr_regfile__rg_mcause [3:0]!=4'd5&& RTL__csr_regfile__rg_mcause [3:0]!=4'd6&& RTL__csr_regfile__rg_mcause [3:0]!=4'd7&& RTL__csr_regfile__rg_mcause [3:0]!=4'd8&& RTL__csr_regfile__rg_mcause [3:0]!=4'd9&& RTL__csr_regfile__rg_mcause [3:0]!=4'd10&& RTL__csr_regfile__rg_mcause [3:0]!=4'd11)$write("unknown interrupt Exc_Code %d", RTL__csr_regfile__rg_mcause [3:0]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd0)$write("INSTRUCTION_ADDR_MISALIGNED");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd1)$write("INSTRUCTION_ACCESS_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd2)$write("ILLEGAL_INSTRUCTION");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd3)$write("BREAKPOINT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd4)$write("LOAD_ADDR_MISALIGNED");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd5)$write("LOAD_ACCESS_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd6)$write("STORE_AMO_ADDR_MISALIGNED");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd7)$write("STORE_AMO_ACCESS_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd8)$write("ECALL_FROM_U");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd9)$write("ECALL_FROM_S");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd11)$write("ECALL_FROM_M");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd12)$write("INSTRUCTION_PAGE_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd13)$write("LOAD_PAGE_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]==4'd15)$write("STORE_AMO_PAGE_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__rg_mcause [4]&& RTL__csr_regfile__rg_mcause [3:0]!=4'd0&& RTL__csr_regfile__rg_mcause [3:0]!=4'd1&& RTL__csr_regfile__rg_mcause [3:0]!=4'd2&& RTL__csr_regfile__rg_mcause [3:0]!=4'd3&& RTL__csr_regfile__rg_mcause [3:0]!=4'd4&& RTL__csr_regfile__rg_mcause [3:0]!=4'd5&& RTL__csr_regfile__rg_mcause [3:0]!=4'd6&& RTL__csr_regfile__rg_mcause [3:0]!=4'd7&& RTL__csr_regfile__rg_mcause [3:0]!=4'd8&& RTL__csr_regfile__rg_mcause [3:0]!=4'd9&& RTL__csr_regfile__rg_mcause [3:0]!=4'd11&& RTL__csr_regfile__rg_mcause [3:0]!=4'd12&& RTL__csr_regfile__rg_mcause [3:0]!=4'd13&& RTL__csr_regfile__rg_mcause [3:0]!=4'd15)$write("unknown trap Exc_Code %d", RTL__csr_regfile__rg_mcause [3:0]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("        ");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" status: 0x%0h", RTL__csr_regfile__csr_mstatus_rg_mstatus );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tvec: 0x%0h",{ RTL__csr_regfile__rg_mtvec [30:1],1'b0, RTL__csr_regfile__rg_mtvec [0]});
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" epc: 0x%0h", RTL__csr_regfile__rg_mepc );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tval: 0x%0h", RTL__csr_regfile__rg_mtval );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("    Return: new pc 0x%0h  ", RTL__csr_regfile__x__h5843 );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" new mstatus:");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("MStatus{","sd:%0d",1'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tsr:%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [22]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tw:%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [21]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tvm:%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [20]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" mxr:%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [19]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" sum:%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [18]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" mprv:%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [17]);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" xs:%0d",2'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" fs:%0d",2'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" mpp:%0d", RTL__csr_regfile__mpp__h7337 );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" spp:%0d",1'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" pies:%0d_%0d%0d", RTL__csr_regfile__csr_mstatus_rg_mstatus [3],1'd0,1'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ies:%0d_%0d%0d",1'd0,1'd0,1'd0);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("}");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" new xcause:");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd0)$write("USER_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd1)$write("SUPERVISOR_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd2)$write("HYPERVISOR_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd3)$write("MACHINE_SW_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd4)$write("USER_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd5)$write("SUPERVISOR_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd6)$write("HYPERVISOR_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd7)$write("MACHINE_TIMER_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd8)$write("USER_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd9)$write("SUPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd10)$write("HYPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL__csr_regfile__csr_trap_actions_nmi && RTL__csr_regfile__csr_trap_actions_interrupt && RTL__csr_regfile__exc_code__h7909 ==4'd11)$write("MACHINE_EXTERNAL_INTERRUPT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__NOT_csr_trap_actions_nmi_97_AND_csr_trap_actio_ETC___d974 )$write("unknown interrupt Exc_Code %d", RTL__csr_regfile__exc_code__h7909 );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd0)$write("INSTRUCTION_ADDR_MISALIGNED");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd1)$write("INSTRUCTION_ACCESS_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd2)$write("ILLEGAL_INSTRUCTION");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd3)$write("BREAKPOINT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd4)$write("LOAD_ADDR_MISALIGNED");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd5)$write("LOAD_ACCESS_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd6)$write("STORE_AMO_ADDR_MISALIGNED");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd7)$write("STORE_AMO_ACCESS_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd8)$write("ECALL_FROM_U");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd9)$write("ECALL_FROM_S");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd11)$write("ECALL_FROM_M");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd12)$write("INSTRUCTION_PAGE_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd13)$write("LOAD_PAGE_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL__csr_regfile__csr_trap_actions_nmi ||! RTL__csr_regfile__csr_trap_actions_interrupt )&& RTL__csr_regfile__exc_code__h7909 ==4'd15)$write("STORE_AMO_PAGE_FAULT");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL__csr_regfile__csr_trap_actions_nmi_OR_NOT_csr_trap_actions_i_ETC___d1025 )$write("unknown trap Exc_Code %d", RTL__csr_regfile__exc_code__h7909 );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" new priv %0d",2'b11);
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_csr_trap_actions && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("");
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__EN_mav_csr_write && RTL__csr_regfile__mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d730 && RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: ERROR: CSR-write addr 0x%0h val 0x%0h not successful", RTL__csr_regfile__rg_mcycle , RTL__csr_regfile__mav_csr_write_csr_addr , RTL__csr_regfile__mav_csr_write_word );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: m_external_interrupt_req: %x", RTL__csr_regfile__rg_mcycle , RTL__csr_regfile__m_external_interrupt_req_set_not_clear );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: s_external_interrupt_req: %x", RTL__csr_regfile__rg_mcycle , RTL__csr_regfile__s_external_interrupt_req_set_not_clear );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: software_interrupt_req: %x", RTL__csr_regfile__rg_mcycle , RTL__csr_regfile__software_interrupt_req_set_not_clear );
             if ( RTL__csr_regfile__RST_N !=1'b0)
                 if ( RTL__csr_regfile__NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: timer_interrupt_req: %x", RTL__csr_regfile__rg_mcycle , RTL__csr_regfile__timer_interrupt_req_set_not_clear );
         end
  assign  RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__rg_state = RTL__csr_regfile__rg_state ; 
  assign  RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__rg_nmi = RTL__csr_regfile__rg_nmi ;
    assign RTL__RTL__DOT__csr_regfile__DOT__rg_nmi = RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__rg_nmi;
    assign RTL__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__csr_regfile__DOT__rg_state = RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__rg_state;
    assign RTL__csr_regfile__CLK = RTL__CLK;
    assign RTL__csr_regfile__RST_N = RTL__RST_N;
    assign RTL__csr_regfile__EN_server_reset_request_put = RTL__csr_regfile$EN_server_reset_request_put;
    assign RTL__csr_regfile$RDY_server_reset_request_put = RTL__csr_regfile__RDY_server_reset_request_put;
    assign RTL__csr_regfile__EN_server_reset_response_get = RTL__csr_regfile$EN_server_reset_response_get;
    assign RTL__csr_regfile$RDY_server_reset_response_get = RTL__csr_regfile__RDY_server_reset_response_get;
    assign RTL__csr_regfile__read_csr_csr_addr = RTL__csr_regfile$read_csr_csr_addr;
    assign RTL__csr_regfile$read_csr = RTL__csr_regfile__read_csr;
    assign RTL__csr_regfile__read_csr_port2_csr_addr = RTL__csr_regfile$read_csr_port2_csr_addr;
    assign RTL__csr_regfile__mav_read_csr_csr_addr = RTL__csr_regfile$mav_read_csr_csr_addr;
    assign RTL__csr_regfile__EN_mav_read_csr = RTL__csr_regfile$EN_mav_read_csr;
    assign RTL__csr_regfile__mav_csr_write_csr_addr = RTL__csr_regfile$mav_csr_write_csr_addr;
    assign RTL__csr_regfile__mav_csr_write_word = RTL__csr_regfile$mav_csr_write_word;
    assign RTL__csr_regfile__EN_mav_csr_write = RTL__csr_regfile$EN_mav_csr_write;
    assign RTL__csr_regfile$read_misa = RTL__csr_regfile__read_misa;
    assign RTL__csr_regfile$read_mstatus = RTL__csr_regfile__read_mstatus;
    assign RTL__csr_regfile$read_satp = RTL__csr_regfile__read_satp;
    assign RTL__csr_regfile__csr_trap_actions_from_priv = RTL__csr_regfile$csr_trap_actions_from_priv;
    assign RTL__csr_regfile__csr_trap_actions_pc = RTL__csr_regfile$csr_trap_actions_pc;
    assign RTL__csr_regfile__csr_trap_actions_nmi = RTL__csr_regfile$csr_trap_actions_nmi;
    assign RTL__csr_regfile__csr_trap_actions_interrupt = RTL__csr_regfile$csr_trap_actions_interrupt;
    assign RTL__csr_regfile__csr_trap_actions_exc_code = RTL__csr_regfile$csr_trap_actions_exc_code;
    assign RTL__csr_regfile__csr_trap_actions_xtval = RTL__csr_regfile$csr_trap_actions_xtval;
    assign RTL__csr_regfile__EN_csr_trap_actions = RTL__csr_regfile$EN_csr_trap_actions;
    assign RTL__csr_regfile$csr_trap_actions = RTL__csr_regfile__csr_trap_actions;
    assign RTL__csr_regfile__csr_ret_actions_from_priv = RTL__csr_regfile$csr_ret_actions_from_priv;
    assign RTL__csr_regfile__EN_csr_ret_actions = RTL__csr_regfile$EN_csr_ret_actions;
    assign RTL__csr_regfile$csr_ret_actions = RTL__csr_regfile__csr_ret_actions;
    assign RTL__csr_regfile$read_csr_minstret = RTL__csr_regfile__read_csr_minstret;
    assign RTL__csr_regfile__EN_csr_minstret_incr = RTL__csr_regfile$EN_csr_minstret_incr;
    assign RTL__csr_regfile$read_csr_mcycle = RTL__csr_regfile__read_csr_mcycle;
    assign RTL__csr_regfile__access_permitted_1_priv = RTL__csr_regfile$access_permitted_1_priv;
    assign RTL__csr_regfile__access_permitted_1_csr_addr = RTL__csr_regfile$access_permitted_1_csr_addr;
    assign RTL__csr_regfile__access_permitted_1_read_not_write = RTL__csr_regfile$access_permitted_1_read_not_write;
    assign RTL__csr_regfile$access_permitted_1 = RTL__csr_regfile__access_permitted_1;
    assign RTL__csr_regfile__access_permitted_2_priv = RTL__csr_regfile$access_permitted_2_priv;
    assign RTL__csr_regfile__access_permitted_2_csr_addr = RTL__csr_regfile$access_permitted_2_csr_addr;
    assign RTL__csr_regfile__access_permitted_2_read_not_write = RTL__csr_regfile$access_permitted_2_read_not_write;
    assign RTL__csr_regfile$access_permitted_2 = RTL__csr_regfile__access_permitted_2;
    assign RTL__csr_regfile__csr_counter_read_fault_priv = RTL__csr_regfile$csr_counter_read_fault_priv;
    assign RTL__csr_regfile__csr_counter_read_fault_csr_addr = RTL__csr_regfile$csr_counter_read_fault_csr_addr;
    assign RTL__csr_regfile__m_external_interrupt_req_set_not_clear = RTL__csr_regfile$m_external_interrupt_req_set_not_clear;
    assign RTL__csr_regfile__s_external_interrupt_req_set_not_clear = RTL__csr_regfile$s_external_interrupt_req_set_not_clear;
    assign RTL__csr_regfile__timer_interrupt_req_set_not_clear = RTL__csr_regfile$timer_interrupt_req_set_not_clear;
    assign RTL__csr_regfile__software_interrupt_req_set_not_clear = RTL__csr_regfile$software_interrupt_req_set_not_clear;
    assign RTL__csr_regfile__interrupt_pending_cur_priv = RTL__csr_regfile$interrupt_pending_cur_priv;
    assign RTL__csr_regfile$interrupt_pending = RTL__csr_regfile__interrupt_pending;
    assign RTL__csr_regfile$wfi_resume = RTL__csr_regfile__wfi_resume;
    assign RTL__csr_regfile__nmi_req_set_not_clear = RTL__csr_regfile$nmi_req_set_not_clear;
    assign RTL__csr_regfile$nmi_pending = RTL__csr_regfile__nmi_pending;
    assign RTL__csr_regfile__EN_debug = RTL__csr_regfile$EN_debug;
      
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;

    parameter RTL__f_reset_reqs__width =1; parameter RTL__f_reset_reqs__guarded =1; 
    reg RTL__f_reset_reqs__full_reg ; 
    reg RTL__f_reset_reqs__empty_reg ; reg[ RTL__f_reset_reqs__width -1:0] RTL__f_reset_reqs__data0_reg ; reg[ RTL__f_reset_reqs__width -1:0] RTL__f_reset_reqs__data1_reg ; 
  assign  RTL__f_reset_reqs__FULL_N = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__EMPTY_N = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__D_OUT = RTL__f_reset_reqs__data0_reg ; 
    wire RTL__f_reset_reqs__d0di =( RTL__f_reset_reqs__ENQ &&! RTL__f_reset_reqs__empty_reg )||( RTL__f_reset_reqs__ENQ && RTL__f_reset_reqs__DEQ && RTL__f_reset_reqs__full_reg ); 
    wire RTL__f_reset_reqs__d0d1 = RTL__f_reset_reqs__DEQ &&! RTL__f_reset_reqs__full_reg ; 
    wire RTL__f_reset_reqs__d0h =((! RTL__f_reset_reqs__DEQ )&&(! RTL__f_reset_reqs__ENQ ))||(! RTL__f_reset_reqs__DEQ && RTL__f_reset_reqs__empty_reg )||(! RTL__f_reset_reqs__ENQ && RTL__f_reset_reqs__full_reg ); 
    wire RTL__f_reset_reqs__d1di = RTL__f_reset_reqs__ENQ & RTL__f_reset_reqs__empty_reg ; 
  always @( posedge  RTL__f_reset_reqs__CLK )
         begin 
             if ( RTL__f_reset_reqs__RST ==1'b0)
                 begin  
                     RTL__f_reset_reqs__empty_reg  <=1'b0; 
                     RTL__f_reset_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__f_reset_reqs__CLR )
                         begin  
                             RTL__f_reset_reqs__empty_reg  <=1'b0; 
                             RTL__f_reset_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__f_reset_reqs__ENQ &&! RTL__f_reset_reqs__DEQ )
                             begin  
                                 RTL__f_reset_reqs__empty_reg  <=1'b1; 
                                 RTL__f_reset_reqs__full_reg  <=! RTL__f_reset_reqs__empty_reg ;
                             end 
                          else 
                             if ( RTL__f_reset_reqs__DEQ &&! RTL__f_reset_reqs__ENQ )
                                 begin  
                                     RTL__f_reset_reqs__full_reg  <=1'b1; 
                                     RTL__f_reset_reqs__empty_reg  <=! RTL__f_reset_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__f_reset_reqs__CLK )
         begin 
             begin  
                 RTL__f_reset_reqs__data0_reg  <={ RTL__f_reset_reqs__width { RTL__f_reset_reqs__d0di }}& RTL__f_reset_reqs__D_IN |{ RTL__f_reset_reqs__width { RTL__f_reset_reqs__d0d1 }}& RTL__f_reset_reqs__data1_reg |{ RTL__f_reset_reqs__width { RTL__f_reset_reqs__d0h }}& RTL__f_reset_reqs__data0_reg ; 
                 RTL__f_reset_reqs__data1_reg  <= RTL__f_reset_reqs__d1di  ?  RTL__f_reset_reqs__D_IN : RTL__f_reset_reqs__data1_reg ;
             end 
         end
  always @( posedge  RTL__f_reset_reqs__CLK )
         begin : RTL__f_reset_reqs__error_checks 
           reg RTL__f_reset_reqs__deqerror , RTL__f_reset_reqs__enqerror ; 
             RTL__f_reset_reqs__deqerror  =0; 
             RTL__f_reset_reqs__enqerror  =0;
             if ( RTL__f_reset_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__f_reset_reqs__empty_reg && RTL__f_reset_reqs__DEQ )
                         begin  
                             RTL__f_reset_reqs__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__f_reset_reqs__full_reg && RTL__f_reset_reqs__ENQ &&(! RTL__f_reset_reqs__DEQ || RTL__f_reset_reqs__guarded ))
                         begin  
                             RTL__f_reset_reqs__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__f_reset_reqs__full_reg ; 
  assign  RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__f_reset_reqs__empty_reg ;
    parameter RTL__f_reset_rsps__width =1; parameter RTL__f_reset_rsps__guarded =1; 
    reg RTL__f_reset_rsps__full_reg ; 
    reg RTL__f_reset_rsps__empty_reg ; reg[ RTL__f_reset_rsps__width -1:0] RTL__f_reset_rsps__data0_reg ; reg[ RTL__f_reset_rsps__width -1:0] RTL__f_reset_rsps__data1_reg ; 
  assign  RTL__f_reset_rsps__FULL_N = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__EMPTY_N = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__D_OUT = RTL__f_reset_rsps__data0_reg ; 
    wire RTL__f_reset_rsps__d0di =( RTL__f_reset_rsps__ENQ &&! RTL__f_reset_rsps__empty_reg )||( RTL__f_reset_rsps__ENQ && RTL__f_reset_rsps__DEQ && RTL__f_reset_rsps__full_reg ); 
    wire RTL__f_reset_rsps__d0d1 = RTL__f_reset_rsps__DEQ &&! RTL__f_reset_rsps__full_reg ; 
    wire RTL__f_reset_rsps__d0h =((! RTL__f_reset_rsps__DEQ )&&(! RTL__f_reset_rsps__ENQ ))||(! RTL__f_reset_rsps__DEQ && RTL__f_reset_rsps__empty_reg )||(! RTL__f_reset_rsps__ENQ && RTL__f_reset_rsps__full_reg ); 
    wire RTL__f_reset_rsps__d1di = RTL__f_reset_rsps__ENQ & RTL__f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__f_reset_rsps__CLK )
         begin 
             if ( RTL__f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__f_reset_rsps__CLR )
                         begin  
                             RTL__f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__f_reset_rsps__ENQ &&! RTL__f_reset_rsps__DEQ )
                             begin  
                                 RTL__f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__f_reset_rsps__full_reg  <=! RTL__f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if ( RTL__f_reset_rsps__DEQ &&! RTL__f_reset_rsps__ENQ )
                                 begin  
                                     RTL__f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__f_reset_rsps__empty_reg  <=! RTL__f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__f_reset_rsps__CLK )
         begin 
             begin  
                 RTL__f_reset_rsps__data0_reg  <={ RTL__f_reset_rsps__width { RTL__f_reset_rsps__d0di }}& RTL__f_reset_rsps__D_IN |{ RTL__f_reset_rsps__width { RTL__f_reset_rsps__d0d1 }}& RTL__f_reset_rsps__data1_reg |{ RTL__f_reset_rsps__width { RTL__f_reset_rsps__d0h }}& RTL__f_reset_rsps__data0_reg ; 
                 RTL__f_reset_rsps__data1_reg  <= RTL__f_reset_rsps__d1di  ?  RTL__f_reset_rsps__D_IN : RTL__f_reset_rsps__data1_reg ;
             end 
         end
  always @( posedge  RTL__f_reset_rsps__CLK )
         begin : RTL__f_reset_rsps__error_checks 
           reg RTL__f_reset_rsps__deqerror , RTL__f_reset_rsps__enqerror ; 
             RTL__f_reset_rsps__deqerror  =0; 
             RTL__f_reset_rsps__enqerror  =0;
             if ( RTL__f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__f_reset_rsps__empty_reg && RTL__f_reset_rsps__DEQ )
                         begin  
                             RTL__f_reset_rsps__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__f_reset_rsps__full_reg && RTL__f_reset_rsps__ENQ &&(! RTL__f_reset_rsps__DEQ || RTL__f_reset_rsps__guarded ))
                         begin  
                             RTL__f_reset_rsps__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__f_reset_rsps__full_reg ; 
  assign  RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__f_reset_rsps__empty_reg ;
    assign RTL__RST_N = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__CLK = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__f_reset_reqs$D_IN = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__f_reset_reqs$ENQ = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__f_reset_reqs$DEQ = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__f_reset_reqs$CLR = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__f_reset_reqs$D_OUT = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__f_reset_reqs$FULL_N = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__f_reset_reqs$EMPTY_N = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__RST_N = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__CLK = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__f_reset_rsps$D_IN = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__f_reset_rsps$ENQ = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__f_reset_rsps$DEQ = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__f_reset_rsps$CLR = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__f_reset_rsps$D_OUT = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__f_reset_rsps$FULL_N = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__f_reset_rsps$EMPTY_N = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
      
    wire RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    wire RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    wire[31:0] RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    wire RTL__gpr_regfile__CLK;
    wire RTL__gpr_regfile__RST_N;
    wire RTL__gpr_regfile__EN_server_reset_request_put;
    wire RTL__gpr_regfile__RDY_server_reset_request_put;
    wire RTL__gpr_regfile__EN_server_reset_response_get;
    wire RTL__gpr_regfile__RDY_server_reset_response_get;
    wire[4:0] RTL__gpr_regfile__read_rs1_rs1;
    wire[31:0] RTL__gpr_regfile__read_rs1;
    wire[4:0] RTL__gpr_regfile__read_rs1_port2_rs1;
    wire[31:0] RTL__gpr_regfile__read_rs1_port2;
    wire[4:0] RTL__gpr_regfile__read_rs2_rs2;
    wire[31:0] RTL__gpr_regfile__read_rs2;
    wire[4:0] RTL__gpr_regfile__write_rd_rd;
    wire[31:0] RTL__gpr_regfile__write_rd_rd_val;
    wire RTL__gpr_regfile__EN_write_rd;

    wire[31:0] RTL__gpr_regfile__read_rs1 , RTL__gpr_regfile__read_rs1_port2 , RTL__gpr_regfile__read_rs2 ; 
    wire RTL__gpr_regfile__RDY_server_reset_request_put , RTL__gpr_regfile__RDY_server_reset_response_get ; reg[1:0] RTL__gpr_regfile__rg_state ; reg[1:0] RTL__gpr_regfile__rg_state$D_IN ; 
    wire RTL__gpr_regfile__rg_state$EN ; 
    wire RTL__gpr_regfile__f_reset_rsps$CLR , RTL__gpr_regfile__f_reset_rsps$DEQ , RTL__gpr_regfile__f_reset_rsps$EMPTY_N , RTL__gpr_regfile__f_reset_rsps$ENQ , RTL__gpr_regfile__f_reset_rsps$FULL_N ; 
    wire[31:0] RTL__gpr_regfile__regfile$D_IN , RTL__gpr_regfile__regfile$D_OUT_1 , RTL__gpr_regfile__regfile$D_OUT_2 , RTL__gpr_regfile__regfile$D_OUT_3 ; 
    wire[4:0] RTL__gpr_regfile__regfile$ADDR_1 , RTL__gpr_regfile__regfile$ADDR_2 , RTL__gpr_regfile__regfile$ADDR_3 , RTL__gpr_regfile__regfile$ADDR_4 , RTL__gpr_regfile__regfile$ADDR_5 , RTL__gpr_regfile__regfile$ADDR_IN ; 
    wire RTL__gpr_regfile__regfile$WE ; 
    wire RTL__gpr_regfile__CAN_FIRE_RL_rl_reset_loop , RTL__gpr_regfile__CAN_FIRE_RL_rl_reset_start , RTL__gpr_regfile__CAN_FIRE_server_reset_request_put , RTL__gpr_regfile__CAN_FIRE_server_reset_response_get , RTL__gpr_regfile__CAN_FIRE_write_rd , RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_loop , RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_start , RTL__gpr_regfile__WILL_FIRE_server_reset_request_put , RTL__gpr_regfile__WILL_FIRE_server_reset_response_get , RTL__gpr_regfile__WILL_FIRE_write_rd ; 
  assign  RTL__gpr_regfile__RDY_server_reset_request_put = RTL__gpr_regfile__f_reset_rsps$FULL_N ; 
  assign  RTL__gpr_regfile__CAN_FIRE_server_reset_request_put = RTL__gpr_regfile__f_reset_rsps$FULL_N ; 
  assign  RTL__gpr_regfile__WILL_FIRE_server_reset_request_put = RTL__gpr_regfile__EN_server_reset_request_put ; 
  assign  RTL__gpr_regfile__RDY_server_reset_response_get = RTL__gpr_regfile__rg_state ==2'd2&& RTL__gpr_regfile__f_reset_rsps$EMPTY_N ; 
  assign  RTL__gpr_regfile__CAN_FIRE_server_reset_response_get = RTL__gpr_regfile__rg_state ==2'd2&& RTL__gpr_regfile__f_reset_rsps$EMPTY_N ; 
  assign  RTL__gpr_regfile__WILL_FIRE_server_reset_response_get = RTL__gpr_regfile__EN_server_reset_response_get ; 
  assign  RTL__gpr_regfile__read_rs1 =( RTL__gpr_regfile__read_rs1_rs1 ==5'd0) ? 32'd0: RTL__gpr_regfile__regfile$D_OUT_3 ; 
  assign  RTL__gpr_regfile__read_rs1_port2 =( RTL__gpr_regfile__read_rs1_port2_rs1 ==5'd0) ? 32'd0: RTL__gpr_regfile__regfile$D_OUT_2 ; 
  assign  RTL__gpr_regfile__read_rs2 =( RTL__gpr_regfile__read_rs2_rs2 ==5'd0) ? 32'd0: RTL__gpr_regfile__regfile$D_OUT_1 ; 
  assign  RTL__gpr_regfile__CAN_FIRE_write_rd =1'd1; 
  assign  RTL__gpr_regfile__WILL_FIRE_write_rd = RTL__gpr_regfile__EN_write_rd ;  
    wire RTL__gpr_regfile__f_reset_rsps__RST;
    wire RTL__gpr_regfile__f_reset_rsps__CLK;
    wire RTL__gpr_regfile__f_reset_rsps__ENQ;
    wire RTL__gpr_regfile__f_reset_rsps__CLR;
    wire RTL__gpr_regfile__f_reset_rsps__DEQ;
    wire RTL__gpr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;

    parameter RTL__gpr_regfile__f_reset_rsps__guarded =1; 
    reg RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
    reg RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__FULL_N = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__EMPTY_N = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__gpr_regfile__f_reset_rsps__CLK )
         begin 
             if ( RTL__gpr_regfile__f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__gpr_regfile__f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__gpr_regfile__f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__gpr_regfile__f_reset_rsps__CLR )
                         begin  
                             RTL__gpr_regfile__f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__gpr_regfile__f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__gpr_regfile__f_reset_rsps__ENQ &&! RTL__gpr_regfile__f_reset_rsps__DEQ )
                             begin  
                                 RTL__gpr_regfile__f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__gpr_regfile__f_reset_rsps__full_reg  <=! RTL__gpr_regfile__f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if (! RTL__gpr_regfile__f_reset_rsps__ENQ && RTL__gpr_regfile__f_reset_rsps__DEQ )
                                 begin  
                                     RTL__gpr_regfile__f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__gpr_regfile__f_reset_rsps__empty_reg  <=! RTL__gpr_regfile__f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__gpr_regfile__f_reset_rsps__CLK )
         begin : RTL__gpr_regfile__f_reset_rsps__error_checks 
           reg RTL__gpr_regfile__f_reset_rsps__deqerror , RTL__gpr_regfile__f_reset_rsps__enqerror ; 
             RTL__gpr_regfile__f_reset_rsps__deqerror  =0; 
             RTL__gpr_regfile__f_reset_rsps__enqerror  =0;
             if ( RTL__gpr_regfile__f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__gpr_regfile__f_reset_rsps__empty_reg && RTL__gpr_regfile__f_reset_rsps__DEQ )
                         begin  
                             RTL__gpr_regfile__f_reset_rsps__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__gpr_regfile__f_reset_rsps__full_reg && RTL__gpr_regfile__f_reset_rsps__ENQ &&(! RTL__gpr_regfile__f_reset_rsps__DEQ || RTL__gpr_regfile__f_reset_rsps__guarded ))
                         begin  
                             RTL__gpr_regfile__f_reset_rsps__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__full_reg ; 
  assign  RTL__gpr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__empty_reg ;
    assign RTL__gpr_regfile__f_reset_rsps__RST = RTL__gpr_regfile__RST_N;
    assign RTL__gpr_regfile__f_reset_rsps__CLK = RTL__gpr_regfile__CLK;
    assign RTL__gpr_regfile__f_reset_rsps__ENQ = RTL__gpr_regfile__f_reset_rsps$ENQ;
    assign RTL__gpr_regfile__f_reset_rsps__CLR = RTL__gpr_regfile__f_reset_rsps$CLR;
    assign RTL__gpr_regfile__f_reset_rsps__DEQ = RTL__gpr_regfile__f_reset_rsps$DEQ;
    assign RTL__gpr_regfile__f_reset_rsps$FULL_N = RTL__gpr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__gpr_regfile__f_reset_rsps$EMPTY_N = RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
      
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    wire[31:0] RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    wire RTL__gpr_regfile__regfile__CLK;
    wire[RTL__gpr_regfile__regfile__addr_width-1:0] RTL__gpr_regfile__regfile__ADDR_IN;
    wire[RTL__gpr_regfile__regfile__data_width-1:0] RTL__gpr_regfile__regfile__D_IN;
    wire RTL__gpr_regfile__regfile__WE;
    wire[RTL__gpr_regfile__regfile__addr_width-1:0] RTL__gpr_regfile__regfile__ADDR_1;
    wire[RTL__gpr_regfile__regfile__data_width-1:0] RTL__gpr_regfile__regfile__D_OUT_1;
    wire[RTL__gpr_regfile__regfile__addr_width-1:0] RTL__gpr_regfile__regfile__ADDR_2;
    wire[RTL__gpr_regfile__regfile__data_width-1:0] RTL__gpr_regfile__regfile__D_OUT_2;
    wire[RTL__gpr_regfile__regfile__addr_width-1:0] RTL__gpr_regfile__regfile__ADDR_3;
    wire[RTL__gpr_regfile__regfile__data_width-1:0] RTL__gpr_regfile__regfile__D_OUT_3;
    wire[RTL__gpr_regfile__regfile__addr_width-1:0] RTL__gpr_regfile__regfile__ADDR_4;
    wire[RTL__gpr_regfile__regfile__data_width-1:0] RTL__gpr_regfile__regfile__D_OUT_4;
    wire[RTL__gpr_regfile__regfile__addr_width-1:0] RTL__gpr_regfile__regfile__ADDR_5;
    wire[RTL__gpr_regfile__regfile__data_width-1:0] RTL__gpr_regfile__regfile__D_OUT_5;

    parameter RTL__gpr_regfile__regfile__addr_width =1; parameter RTL__gpr_regfile__regfile__data_width =1; parameter RTL__gpr_regfile__regfile__lo =0; parameter RTL__gpr_regfile__regfile__hi =1; reg[ RTL__gpr_regfile__regfile__data_width -1:0] RTL__gpr_regfile__regfile__arr [ RTL__gpr_regfile__regfile__lo : RTL__gpr_regfile__regfile__hi ]; 
  always @( posedge  RTL__gpr_regfile__regfile__CLK )
         begin 
             if ( RTL__gpr_regfile__regfile__WE ) 
                 RTL__gpr_regfile__regfile__arr  [ RTL__gpr_regfile__regfile__ADDR_IN ]<= RTL__gpr_regfile__regfile__D_IN ;
         end
  assign  RTL__gpr_regfile__regfile__D_OUT_1 = RTL__gpr_regfile__regfile__arr [ RTL__gpr_regfile__regfile__ADDR_1 ]; 
  assign  RTL__gpr_regfile__regfile__D_OUT_2 = RTL__gpr_regfile__regfile__arr [ RTL__gpr_regfile__regfile__ADDR_2 ]; 
  assign  RTL__gpr_regfile__regfile__D_OUT_3 = RTL__gpr_regfile__regfile__arr [ RTL__gpr_regfile__regfile__ADDR_3 ]; 
  assign  RTL__gpr_regfile__regfile__D_OUT_4 = RTL__gpr_regfile__regfile__arr [ RTL__gpr_regfile__regfile__ADDR_4 ]; 
  assign  RTL__gpr_regfile__regfile__D_OUT_5 = RTL__gpr_regfile__regfile__arr [ RTL__gpr_regfile__regfile__ADDR_5 ]; 
  always @( posedge  RTL__gpr_regfile__regfile__CLK )
         begin : RTL__gpr_regfile__regfile__runtime_check 
           reg RTL__gpr_regfile__regfile__enable_check ; 
             RTL__gpr_regfile__regfile__enable_check  =0;
             if ( RTL__gpr_regfile__regfile__enable_check )
                 begin 
                     if (( RTL__gpr_regfile__regfile__ADDR_1 < RTL__gpr_regfile__regfile__lo )||( RTL__gpr_regfile__regfile__ADDR_1 > RTL__gpr_regfile__regfile__hi ))$display("Warning: RegFile: %m -- Address port 1 is out of bounds: %h", RTL__gpr_regfile__regfile__ADDR_1 );
                     if (( RTL__gpr_regfile__regfile__ADDR_2 < RTL__gpr_regfile__regfile__lo )||( RTL__gpr_regfile__regfile__ADDR_2 > RTL__gpr_regfile__regfile__hi ))$display("Warning: RegFile: %m -- Address port 2 is out of bounds: %h", RTL__gpr_regfile__regfile__ADDR_2 );
                     if (( RTL__gpr_regfile__regfile__ADDR_3 < RTL__gpr_regfile__regfile__lo )||( RTL__gpr_regfile__regfile__ADDR_3 > RTL__gpr_regfile__regfile__hi ))$display("Warning: RegFile: %m -- Address port 3 is out of bounds: %h", RTL__gpr_regfile__regfile__ADDR_3 );
                     if (( RTL__gpr_regfile__regfile__ADDR_4 < RTL__gpr_regfile__regfile__lo )||( RTL__gpr_regfile__regfile__ADDR_4 > RTL__gpr_regfile__regfile__hi ))$display("Warning: RegFile: %m -- Address port 4 is out of bounds: %h", RTL__gpr_regfile__regfile__ADDR_4 );
                     if (( RTL__gpr_regfile__regfile__ADDR_5 < RTL__gpr_regfile__regfile__lo )||( RTL__gpr_regfile__regfile__ADDR_5 > RTL__gpr_regfile__regfile__hi ))$display("Warning: RegFile: %m -- Address port 5 is out of bounds: %h", RTL__gpr_regfile__regfile__ADDR_5 );
                     if ( RTL__gpr_regfile__regfile__WE &&( RTL__gpr_regfile__regfile__ADDR_IN < RTL__gpr_regfile__regfile__lo )||( RTL__gpr_regfile__regfile__ADDR_IN > RTL__gpr_regfile__regfile__hi ))$display("Warning: RegFile: %m -- Write Address port is out of bounds: %h", RTL__gpr_regfile__regfile__ADDR_IN );
                 end 
         end
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL__gpr_regfile__regfile__arr [15]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL__gpr_regfile__regfile__arr [12]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL__gpr_regfile__regfile__arr [7]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL__gpr_regfile__regfile__arr [10]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL__gpr_regfile__regfile__arr [1]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL__gpr_regfile__regfile__arr [6]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL__gpr_regfile__regfile__arr [31]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL__gpr_regfile__regfile__arr [29]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL__gpr_regfile__regfile__arr [27]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL__gpr_regfile__regfile__arr [25]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL__gpr_regfile__regfile__arr [23]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL__gpr_regfile__regfile__arr [22]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL__gpr_regfile__regfile__arr [21]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL__gpr_regfile__regfile__arr [18]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL__gpr_regfile__regfile__arr [16]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL__gpr_regfile__regfile__arr [28]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL__gpr_regfile__regfile__arr [2]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL__gpr_regfile__regfile__arr [24]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL__gpr_regfile__regfile__arr [30]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL__gpr_regfile__regfile__arr [26]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL__gpr_regfile__regfile__arr [13]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL__gpr_regfile__regfile__arr [19]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL__gpr_regfile__regfile__arr [5]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL__gpr_regfile__regfile__arr [20]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL__gpr_regfile__regfile__arr [4]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL__gpr_regfile__regfile__arr [11]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL__gpr_regfile__regfile__arr [8]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL__gpr_regfile__regfile__arr [3]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL__gpr_regfile__regfile__arr [9]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL__gpr_regfile__regfile__arr [14]; 
  assign  RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL__gpr_regfile__regfile__arr [17];
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    assign RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL__gpr_regfile__regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    assign RTL__gpr_regfile__regfile__CLK = RTL__gpr_regfile__CLK;
    assign RTL__gpr_regfile__regfile__ADDR_IN = RTL__gpr_regfile__regfile$ADDR_IN;
    assign RTL__gpr_regfile__regfile__D_IN = RTL__gpr_regfile__regfile$D_IN;
    assign RTL__gpr_regfile__regfile__WE = RTL__gpr_regfile__regfile$WE;
    assign RTL__gpr_regfile__regfile__ADDR_1 = RTL__gpr_regfile__regfile$ADDR_1;
    assign RTL__gpr_regfile__regfile$D_OUT_1 = RTL__gpr_regfile__regfile__D_OUT_1;
    assign RTL__gpr_regfile__regfile__ADDR_2 = RTL__gpr_regfile__regfile$ADDR_2;
    assign RTL__gpr_regfile__regfile$D_OUT_2 = RTL__gpr_regfile__regfile__D_OUT_2;
    assign RTL__gpr_regfile__regfile__ADDR_3 = RTL__gpr_regfile__regfile$ADDR_3;
    assign RTL__gpr_regfile__regfile$D_OUT_3 = RTL__gpr_regfile__regfile__D_OUT_3;
    assign RTL__gpr_regfile__regfile__ADDR_4 = RTL__gpr_regfile__regfile$ADDR_4;
    assign RTL__gpr_regfile__regfile__ADDR_5 = RTL__gpr_regfile__regfile$ADDR_5;
     
  assign  RTL__gpr_regfile__CAN_FIRE_RL_rl_reset_start = RTL__gpr_regfile__rg_state ==2'd0; 
  assign  RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_start = RTL__gpr_regfile__rg_state ==2'd0; 
  assign  RTL__gpr_regfile__CAN_FIRE_RL_rl_reset_loop = RTL__gpr_regfile__rg_state ==2'd1; 
  assign  RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_loop = RTL__gpr_regfile__rg_state ==2'd1; 
  always @(    RTL__gpr_regfile__EN_server_reset_request_put              or   RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_loop           or   RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_start  )
         case (1'b1) 
          RTL__gpr_regfile__EN_server_reset_request_put  : 
              RTL__gpr_regfile__rg_state$D_IN  =2'd0; 
          RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_loop  : 
              RTL__gpr_regfile__rg_state$D_IN  =2'd2; 
          RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_start  : 
              RTL__gpr_regfile__rg_state$D_IN  =2'd1;
          default : 
              RTL__gpr_regfile__rg_state$D_IN  =2'b10;endcase
  assign  RTL__gpr_regfile__rg_state$EN = RTL__gpr_regfile__EN_server_reset_request_put || RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_start || RTL__gpr_regfile__WILL_FIRE_RL_rl_reset_loop ; 
  assign  RTL__gpr_regfile__f_reset_rsps$ENQ = RTL__gpr_regfile__EN_server_reset_request_put ; 
  assign  RTL__gpr_regfile__f_reset_rsps$DEQ = RTL__gpr_regfile__EN_server_reset_response_get ; 
  assign  RTL__gpr_regfile__f_reset_rsps$CLR =1'b0; 
  assign  RTL__gpr_regfile__regfile$ADDR_1 = RTL__gpr_regfile__read_rs2_rs2 ; 
  assign  RTL__gpr_regfile__regfile$ADDR_2 = RTL__gpr_regfile__read_rs1_port2_rs1 ; 
  assign  RTL__gpr_regfile__regfile$ADDR_3 = RTL__gpr_regfile__read_rs1_rs1 ; 
  assign  RTL__gpr_regfile__regfile$ADDR_4 =5'h0; 
  assign  RTL__gpr_regfile__regfile$ADDR_5 =5'h0; 
  assign  RTL__gpr_regfile__regfile$ADDR_IN = RTL__gpr_regfile__write_rd_rd ; 
  assign  RTL__gpr_regfile__regfile$D_IN = RTL__gpr_regfile__write_rd_rd_val ; 
  assign  RTL__gpr_regfile__regfile$WE = RTL__gpr_regfile__EN_write_rd && RTL__gpr_regfile__write_rd_rd !=5'd0; 
  always @( posedge  RTL__gpr_regfile__CLK )
         begin 
             if ( RTL__gpr_regfile__RST_N ==1'b0)
                 begin  
                     RTL__gpr_regfile__rg_state  <=2'd0;
                 end 
              else 
                 begin 
                     if ( RTL__gpr_regfile__rg_state$EN ) 
                         RTL__gpr_regfile__rg_state  <= RTL__gpr_regfile__rg_state$D_IN ;
                 end 
         end
 
    assign RTL__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    assign RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL__gpr_regfile__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    assign RTL__gpr_regfile__CLK = RTL__CLK;
    assign RTL__gpr_regfile__RST_N = RTL__RST_N;
    assign RTL__gpr_regfile__EN_server_reset_request_put = RTL__gpr_regfile$EN_server_reset_request_put;
    assign RTL__gpr_regfile$RDY_server_reset_request_put = RTL__gpr_regfile__RDY_server_reset_request_put;
    assign RTL__gpr_regfile__EN_server_reset_response_get = RTL__gpr_regfile$EN_server_reset_response_get;
    assign RTL__gpr_regfile$RDY_server_reset_response_get = RTL__gpr_regfile__RDY_server_reset_response_get;
    assign RTL__gpr_regfile__read_rs1_rs1 = RTL__gpr_regfile$read_rs1_rs1;
    assign RTL__gpr_regfile$read_rs1 = RTL__gpr_regfile__read_rs1;
    assign RTL__gpr_regfile__read_rs1_port2_rs1 = RTL__gpr_regfile$read_rs1_port2_rs1;
    assign RTL__gpr_regfile__read_rs2_rs2 = RTL__gpr_regfile$read_rs2_rs2;
    assign RTL__gpr_regfile$read_rs2 = RTL__gpr_regfile__read_rs2;
    assign RTL__gpr_regfile__write_rd_rd = RTL__gpr_regfile$write_rd_rd;
    assign RTL__gpr_regfile__write_rd_rd_val = RTL__gpr_regfile$write_rd_rd_val;
    assign RTL__gpr_regfile__EN_write_rd = RTL__gpr_regfile$EN_write_rd;
      
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire[31:0] RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire[31:0] RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__CLK;
    wire RTL__near_mem__RST_N;
    wire RTL__near_mem__EN_server_reset_request_put;
    wire RTL__near_mem__RDY_server_reset_request_put;
    wire RTL__near_mem__EN_server_reset_response_get;
    wire RTL__near_mem__RDY_server_reset_response_get;
    wire[2:0] RTL__near_mem__imem_req_f3;
    wire[31:0] RTL__near_mem__imem_req_addr;
    wire[1:0] RTL__near_mem__imem_req_priv;
    wire RTL__near_mem__imem_req_sstatus_SUM;
    wire RTL__near_mem__imem_req_mstatus_MXR;
    wire[31:0] RTL__near_mem__imem_req_satp;
    wire RTL__near_mem__EN_imem_req;
    wire RTL__near_mem__imem_valid;
    wire RTL__near_mem__imem_is_i32_not_i16;
    wire[31:0] RTL__near_mem__imem_pc;
    wire[31:0] RTL__near_mem__imem_instr;
    wire RTL__near_mem__imem_exc;
    wire[3:0] RTL__near_mem__imem_exc_code;
    wire[31:0] RTL__near_mem__imem_tval;
    wire RTL__near_mem__imem_master_awvalid;
    wire[3:0] RTL__near_mem__imem_master_awid;
    wire[63:0] RTL__near_mem__imem_master_awaddr;
    wire[7:0] RTL__near_mem__imem_master_awlen;
    wire[2:0] RTL__near_mem__imem_master_awsize;
    wire[1:0] RTL__near_mem__imem_master_awburst;
    wire RTL__near_mem__imem_master_awlock;
    wire[3:0] RTL__near_mem__imem_master_awcache;
    wire[2:0] RTL__near_mem__imem_master_awprot;
    wire[3:0] RTL__near_mem__imem_master_awqos;
    wire[3:0] RTL__near_mem__imem_master_awregion;
    wire RTL__near_mem__imem_master_awready;
    wire RTL__near_mem__imem_master_wvalid;
    wire[63:0] RTL__near_mem__imem_master_wdata;
    wire[7:0] RTL__near_mem__imem_master_wstrb;
    wire RTL__near_mem__imem_master_wlast;
    wire RTL__near_mem__imem_master_wready;
    wire RTL__near_mem__imem_master_bvalid;
    wire[3:0] RTL__near_mem__imem_master_bid;
    wire[1:0] RTL__near_mem__imem_master_bresp;
    wire RTL__near_mem__imem_master_bready;
    wire RTL__near_mem__imem_master_arvalid;
    wire[3:0] RTL__near_mem__imem_master_arid;
    wire[63:0] RTL__near_mem__imem_master_araddr;
    wire[7:0] RTL__near_mem__imem_master_arlen;
    wire[2:0] RTL__near_mem__imem_master_arsize;
    wire[1:0] RTL__near_mem__imem_master_arburst;
    wire RTL__near_mem__imem_master_arlock;
    wire[3:0] RTL__near_mem__imem_master_arcache;
    wire[2:0] RTL__near_mem__imem_master_arprot;
    wire[3:0] RTL__near_mem__imem_master_arqos;
    wire[3:0] RTL__near_mem__imem_master_arregion;
    wire RTL__near_mem__imem_master_arready;
    wire RTL__near_mem__imem_master_rvalid;
    wire[3:0] RTL__near_mem__imem_master_rid;
    wire[63:0] RTL__near_mem__imem_master_rdata;
    wire[1:0] RTL__near_mem__imem_master_rresp;
    wire RTL__near_mem__imem_master_rlast;
    wire RTL__near_mem__imem_master_rready;
    wire RTL__near_mem__dmem_req_op;
    wire[2:0] RTL__near_mem__dmem_req_f3;
    wire[31:0] RTL__near_mem__dmem_req_addr;
    wire[63:0] RTL__near_mem__dmem_req_store_value;
    wire[1:0] RTL__near_mem__dmem_req_priv;
    wire RTL__near_mem__dmem_req_sstatus_SUM;
    wire RTL__near_mem__dmem_req_mstatus_MXR;
    wire[31:0] RTL__near_mem__dmem_req_satp;
    wire RTL__near_mem__EN_dmem_req;
    wire RTL__near_mem__dmem_valid;
    wire[63:0] RTL__near_mem__dmem_word64;
    wire[63:0] RTL__near_mem__dmem_st_amo_val;
    wire RTL__near_mem__dmem_exc;
    wire[3:0] RTL__near_mem__dmem_exc_code;
    wire RTL__near_mem__dmem_master_awvalid;
    wire[3:0] RTL__near_mem__dmem_master_awid;
    wire[63:0] RTL__near_mem__dmem_master_awaddr;
    wire[7:0] RTL__near_mem__dmem_master_awlen;
    wire[2:0] RTL__near_mem__dmem_master_awsize;
    wire[1:0] RTL__near_mem__dmem_master_awburst;
    wire RTL__near_mem__dmem_master_awlock;
    wire[3:0] RTL__near_mem__dmem_master_awcache;
    wire[2:0] RTL__near_mem__dmem_master_awprot;
    wire[3:0] RTL__near_mem__dmem_master_awqos;
    wire[3:0] RTL__near_mem__dmem_master_awregion;
    wire RTL__near_mem__dmem_master_awready;
    wire RTL__near_mem__dmem_master_wvalid;
    wire[63:0] RTL__near_mem__dmem_master_wdata;
    wire[7:0] RTL__near_mem__dmem_master_wstrb;
    wire RTL__near_mem__dmem_master_wlast;
    wire RTL__near_mem__dmem_master_wready;
    wire RTL__near_mem__dmem_master_bvalid;
    wire[3:0] RTL__near_mem__dmem_master_bid;
    wire[1:0] RTL__near_mem__dmem_master_bresp;
    wire RTL__near_mem__dmem_master_bready;
    wire RTL__near_mem__dmem_master_arvalid;
    wire[3:0] RTL__near_mem__dmem_master_arid;
    wire[63:0] RTL__near_mem__dmem_master_araddr;
    wire[7:0] RTL__near_mem__dmem_master_arlen;
    wire[2:0] RTL__near_mem__dmem_master_arsize;
    wire[1:0] RTL__near_mem__dmem_master_arburst;
    wire RTL__near_mem__dmem_master_arlock;
    wire[3:0] RTL__near_mem__dmem_master_arcache;
    wire[2:0] RTL__near_mem__dmem_master_arprot;
    wire[3:0] RTL__near_mem__dmem_master_arqos;
    wire[3:0] RTL__near_mem__dmem_master_arregion;
    wire RTL__near_mem__dmem_master_arready;
    wire RTL__near_mem__dmem_master_rvalid;
    wire[3:0] RTL__near_mem__dmem_master_rid;
    wire[63:0] RTL__near_mem__dmem_master_rdata;
    wire[1:0] RTL__near_mem__dmem_master_rresp;
    wire RTL__near_mem__dmem_master_rlast;
    wire RTL__near_mem__dmem_master_rready;
    wire RTL__near_mem__EN_server_fence_i_request_put;
    wire RTL__near_mem__RDY_server_fence_i_request_put;
    wire RTL__near_mem__EN_server_fence_i_response_get;
    wire RTL__near_mem__RDY_server_fence_i_response_get;
    wire[7:0] RTL__near_mem__server_fence_request_put;
    wire RTL__near_mem__EN_server_fence_request_put;
    wire RTL__near_mem__RDY_server_fence_request_put;
    wire RTL__near_mem__EN_server_fence_response_get;
    wire RTL__near_mem__RDY_server_fence_response_get;
    wire RTL__near_mem__EN_sfence_vma;
    wire RTL__near_mem__RDY_sfence_vma;

    wire[63:0] RTL__near_mem__dmem_master_araddr , RTL__near_mem__dmem_master_awaddr , RTL__near_mem__dmem_master_wdata , RTL__near_mem__dmem_st_amo_val , RTL__near_mem__dmem_word64 , RTL__near_mem__imem_master_araddr , RTL__near_mem__imem_master_awaddr , RTL__near_mem__imem_master_wdata ; 
    wire[31:0] RTL__near_mem__imem_instr , RTL__near_mem__imem_pc , RTL__near_mem__imem_tval ; 
    wire[7:0] RTL__near_mem__dmem_master_arlen , RTL__near_mem__dmem_master_awlen , RTL__near_mem__dmem_master_wstrb , RTL__near_mem__imem_master_arlen , RTL__near_mem__imem_master_awlen , RTL__near_mem__imem_master_wstrb ; 
    wire[3:0] RTL__near_mem__dmem_exc_code , RTL__near_mem__dmem_master_arcache , RTL__near_mem__dmem_master_arid , RTL__near_mem__dmem_master_arqos , RTL__near_mem__dmem_master_arregion , RTL__near_mem__dmem_master_awcache , RTL__near_mem__dmem_master_awid , RTL__near_mem__dmem_master_awqos , RTL__near_mem__dmem_master_awregion , RTL__near_mem__imem_exc_code , RTL__near_mem__imem_master_arcache , RTL__near_mem__imem_master_arid , RTL__near_mem__imem_master_arqos , RTL__near_mem__imem_master_arregion , RTL__near_mem__imem_master_awcache , RTL__near_mem__imem_master_awid , RTL__near_mem__imem_master_awqos , RTL__near_mem__imem_master_awregion ; 
    wire[2:0] RTL__near_mem__dmem_master_arprot , RTL__near_mem__dmem_master_arsize , RTL__near_mem__dmem_master_awprot , RTL__near_mem__dmem_master_awsize , RTL__near_mem__imem_master_arprot , RTL__near_mem__imem_master_arsize , RTL__near_mem__imem_master_awprot , RTL__near_mem__imem_master_awsize ; 
    wire[1:0] RTL__near_mem__dmem_master_arburst , RTL__near_mem__dmem_master_awburst , RTL__near_mem__imem_master_arburst , RTL__near_mem__imem_master_awburst ; 
    wire RTL__near_mem__RDY_server_fence_i_request_put , RTL__near_mem__RDY_server_fence_i_response_get , RTL__near_mem__RDY_server_fence_request_put , RTL__near_mem__RDY_server_fence_response_get , RTL__near_mem__RDY_server_reset_request_put , RTL__near_mem__RDY_server_reset_response_get , RTL__near_mem__RDY_sfence_vma , RTL__near_mem__dmem_exc , RTL__near_mem__dmem_master_arlock , RTL__near_mem__dmem_master_arvalid , RTL__near_mem__dmem_master_awlock , RTL__near_mem__dmem_master_awvalid , RTL__near_mem__dmem_master_bready , RTL__near_mem__dmem_master_rready , RTL__near_mem__dmem_master_wlast , RTL__near_mem__dmem_master_wvalid , RTL__near_mem__dmem_valid , RTL__near_mem__imem_exc , RTL__near_mem__imem_is_i32_not_i16 , RTL__near_mem__imem_master_arlock , RTL__near_mem__imem_master_arvalid , RTL__near_mem__imem_master_awlock , RTL__near_mem__imem_master_awvalid , RTL__near_mem__imem_master_bready , RTL__near_mem__imem_master_rready , RTL__near_mem__imem_master_wlast , RTL__near_mem__imem_master_wvalid , RTL__near_mem__imem_valid ; reg[3:0] RTL__near_mem__cfg_verbosity ; 
    wire[3:0] RTL__near_mem__cfg_verbosity$D_IN ; 
    wire RTL__near_mem__cfg_verbosity$EN ; reg[1:0] RTL__near_mem__rg_state ; reg[1:0] RTL__near_mem__rg_state$D_IN ; 
    wire RTL__near_mem__rg_state$EN ; 
    wire[63:0] RTL__near_mem__dcache$mem_master_araddr , RTL__near_mem__dcache$mem_master_awaddr , RTL__near_mem__dcache$mem_master_rdata , RTL__near_mem__dcache$mem_master_wdata , RTL__near_mem__dcache$req_st_value , RTL__near_mem__dcache$word64 ; 
    wire[31:0] RTL__near_mem__dcache$req_addr , RTL__near_mem__dcache$req_satp ; 
    wire[7:0] RTL__near_mem__dcache$mem_master_arlen , RTL__near_mem__dcache$mem_master_awlen , RTL__near_mem__dcache$mem_master_wstrb ; 
    wire[3:0] RTL__near_mem__dcache$exc_code , RTL__near_mem__dcache$mem_master_arcache , RTL__near_mem__dcache$mem_master_arid , RTL__near_mem__dcache$mem_master_arqos , RTL__near_mem__dcache$mem_master_arregion , RTL__near_mem__dcache$mem_master_awcache , RTL__near_mem__dcache$mem_master_awid , RTL__near_mem__dcache$mem_master_awqos , RTL__near_mem__dcache$mem_master_awregion , RTL__near_mem__dcache$mem_master_bid , RTL__near_mem__dcache$mem_master_rid , RTL__near_mem__dcache$set_verbosity_verbosity ; 
    wire[2:0] RTL__near_mem__dcache$mem_master_arprot , RTL__near_mem__dcache$mem_master_arsize , RTL__near_mem__dcache$mem_master_awprot , RTL__near_mem__dcache$mem_master_awsize , RTL__near_mem__dcache$req_f3 ; 
    wire[1:0] RTL__near_mem__dcache$mem_master_arburst , RTL__near_mem__dcache$mem_master_awburst , RTL__near_mem__dcache$mem_master_bresp , RTL__near_mem__dcache$mem_master_rresp , RTL__near_mem__dcache$req_priv ; 
    wire RTL__near_mem__dcache$EN_req , RTL__near_mem__dcache$EN_server_flush_request_put , RTL__near_mem__dcache$EN_server_flush_response_get , RTL__near_mem__dcache$EN_server_reset_request_put , RTL__near_mem__dcache$EN_server_reset_response_get , RTL__near_mem__dcache$EN_set_verbosity , RTL__near_mem__dcache$EN_tlb_flush , RTL__near_mem__dcache$RDY_server_flush_request_put , RTL__near_mem__dcache$RDY_server_flush_response_get , RTL__near_mem__dcache$RDY_server_reset_request_put , RTL__near_mem__dcache$RDY_server_reset_response_get , RTL__near_mem__dcache$exc , RTL__near_mem__dcache$mem_master_arlock , RTL__near_mem__dcache$mem_master_arready , RTL__near_mem__dcache$mem_master_arvalid , RTL__near_mem__dcache$mem_master_awlock , RTL__near_mem__dcache$mem_master_awready , RTL__near_mem__dcache$mem_master_awvalid , RTL__near_mem__dcache$mem_master_bready , RTL__near_mem__dcache$mem_master_bvalid , RTL__near_mem__dcache$mem_master_rlast , RTL__near_mem__dcache$mem_master_rready , RTL__near_mem__dcache$mem_master_rvalid , RTL__near_mem__dcache$mem_master_wlast , RTL__near_mem__dcache$mem_master_wready , RTL__near_mem__dcache$mem_master_wvalid , RTL__near_mem__dcache$req_mstatus_MXR , RTL__near_mem__dcache$req_op , RTL__near_mem__dcache$req_sstatus_SUM , RTL__near_mem__dcache$valid ; 
    wire RTL__near_mem__f_reset_rsps$CLR , RTL__near_mem__f_reset_rsps$DEQ , RTL__near_mem__f_reset_rsps$EMPTY_N , RTL__near_mem__f_reset_rsps$ENQ , RTL__near_mem__f_reset_rsps$FULL_N ; 
    wire[63:0] RTL__near_mem__icache$mem_master_araddr , RTL__near_mem__icache$mem_master_awaddr , RTL__near_mem__icache$mem_master_rdata , RTL__near_mem__icache$mem_master_wdata , RTL__near_mem__icache$req_st_value , RTL__near_mem__icache$word64 ; 
    wire[31:0] RTL__near_mem__icache$addr , RTL__near_mem__icache$req_addr , RTL__near_mem__icache$req_satp ; 
    wire[7:0] RTL__near_mem__icache$mem_master_arlen , RTL__near_mem__icache$mem_master_awlen , RTL__near_mem__icache$mem_master_wstrb ; 
    wire[3:0] RTL__near_mem__icache$exc_code , RTL__near_mem__icache$mem_master_arcache , RTL__near_mem__icache$mem_master_arid , RTL__near_mem__icache$mem_master_arqos , RTL__near_mem__icache$mem_master_arregion , RTL__near_mem__icache$mem_master_awcache , RTL__near_mem__icache$mem_master_awid , RTL__near_mem__icache$mem_master_awqos , RTL__near_mem__icache$mem_master_awregion , RTL__near_mem__icache$mem_master_bid , RTL__near_mem__icache$mem_master_rid , RTL__near_mem__icache$set_verbosity_verbosity ; 
    wire[2:0] RTL__near_mem__icache$mem_master_arprot , RTL__near_mem__icache$mem_master_arsize , RTL__near_mem__icache$mem_master_awprot , RTL__near_mem__icache$mem_master_awsize , RTL__near_mem__icache$req_f3 ; 
    wire[1:0] RTL__near_mem__icache$mem_master_arburst , RTL__near_mem__icache$mem_master_awburst , RTL__near_mem__icache$mem_master_bresp , RTL__near_mem__icache$mem_master_rresp , RTL__near_mem__icache$req_priv ; 
    wire RTL__near_mem__icache$EN_req , RTL__near_mem__icache$EN_server_flush_request_put , RTL__near_mem__icache$EN_server_flush_response_get , RTL__near_mem__icache$EN_server_reset_request_put , RTL__near_mem__icache$EN_server_reset_response_get , RTL__near_mem__icache$EN_set_verbosity , RTL__near_mem__icache$EN_tlb_flush , RTL__near_mem__icache$RDY_server_flush_request_put , RTL__near_mem__icache$RDY_server_flush_response_get , RTL__near_mem__icache$RDY_server_reset_request_put , RTL__near_mem__icache$RDY_server_reset_response_get , RTL__near_mem__icache$exc , RTL__near_mem__icache$mem_master_arlock , RTL__near_mem__icache$mem_master_arready , RTL__near_mem__icache$mem_master_arvalid , RTL__near_mem__icache$mem_master_awlock , RTL__near_mem__icache$mem_master_awready , RTL__near_mem__icache$mem_master_awvalid , RTL__near_mem__icache$mem_master_bready , RTL__near_mem__icache$mem_master_bvalid , RTL__near_mem__icache$mem_master_rlast , RTL__near_mem__icache$mem_master_rready , RTL__near_mem__icache$mem_master_rvalid , RTL__near_mem__icache$mem_master_wlast , RTL__near_mem__icache$mem_master_wready , RTL__near_mem__icache$mem_master_wvalid , RTL__near_mem__icache$req_mstatus_MXR , RTL__near_mem__icache$req_op , RTL__near_mem__icache$req_sstatus_SUM , RTL__near_mem__icache$valid ; 
    wire[63:0] RTL__near_mem__soc_map$m_is_IO_addr_addr , RTL__near_mem__soc_map$m_is_mem_addr_addr , RTL__near_mem__soc_map$m_is_near_mem_IO_addr_addr ; 
    wire RTL__near_mem__CAN_FIRE_RL_rl_reset , RTL__near_mem__CAN_FIRE_RL_rl_reset_complete , RTL__near_mem__CAN_FIRE_dmem_master_m_arready , RTL__near_mem__CAN_FIRE_dmem_master_m_awready , RTL__near_mem__CAN_FIRE_dmem_master_m_bvalid , RTL__near_mem__CAN_FIRE_dmem_master_m_rvalid , RTL__near_mem__CAN_FIRE_dmem_master_m_wready , RTL__near_mem__CAN_FIRE_dmem_req , RTL__near_mem__CAN_FIRE_imem_master_m_arready , RTL__near_mem__CAN_FIRE_imem_master_m_awready , RTL__near_mem__CAN_FIRE_imem_master_m_bvalid , RTL__near_mem__CAN_FIRE_imem_master_m_rvalid , RTL__near_mem__CAN_FIRE_imem_master_m_wready , RTL__near_mem__CAN_FIRE_imem_req , RTL__near_mem__CAN_FIRE_server_fence_i_request_put , RTL__near_mem__CAN_FIRE_server_fence_i_response_get , RTL__near_mem__CAN_FIRE_server_fence_request_put , RTL__near_mem__CAN_FIRE_server_fence_response_get , RTL__near_mem__CAN_FIRE_server_reset_request_put , RTL__near_mem__CAN_FIRE_server_reset_response_get , RTL__near_mem__CAN_FIRE_sfence_vma , RTL__near_mem__WILL_FIRE_RL_rl_reset , RTL__near_mem__WILL_FIRE_RL_rl_reset_complete , RTL__near_mem__WILL_FIRE_dmem_master_m_arready , RTL__near_mem__WILL_FIRE_dmem_master_m_awready , RTL__near_mem__WILL_FIRE_dmem_master_m_bvalid , RTL__near_mem__WILL_FIRE_dmem_master_m_rvalid , RTL__near_mem__WILL_FIRE_dmem_master_m_wready , RTL__near_mem__WILL_FIRE_dmem_req , RTL__near_mem__WILL_FIRE_imem_master_m_arready , RTL__near_mem__WILL_FIRE_imem_master_m_awready , RTL__near_mem__WILL_FIRE_imem_master_m_bvalid , RTL__near_mem__WILL_FIRE_imem_master_m_rvalid , RTL__near_mem__WILL_FIRE_imem_master_m_wready , RTL__near_mem__WILL_FIRE_imem_req , RTL__near_mem__WILL_FIRE_server_fence_i_request_put , RTL__near_mem__WILL_FIRE_server_fence_i_response_get , RTL__near_mem__WILL_FIRE_server_fence_request_put , RTL__near_mem__WILL_FIRE_server_fence_response_get , RTL__near_mem__WILL_FIRE_server_reset_request_put , RTL__near_mem__WILL_FIRE_server_reset_response_get , RTL__near_mem__WILL_FIRE_sfence_vma ; 
    wire RTL__near_mem__MUX_rg_state$write_1__SEL_2 , RTL__near_mem__MUX_rg_state$write_1__SEL_3 ; reg[31:0] RTL__near_mem__v__h1643 ; reg[31:0] RTL__near_mem__v__h1794 ; reg[31:0] RTL__near_mem__v__h1637 ; reg[31:0] RTL__near_mem__v__h1788 ; 
    wire RTL__near_mem__NOT_cfg_verbosity_read_ULE_1___d9 ; 
  assign  RTL__near_mem__RDY_server_reset_request_put = RTL__near_mem__rg_state ==2'd2; 
  assign  RTL__near_mem__CAN_FIRE_server_reset_request_put = RTL__near_mem__rg_state ==2'd2; 
  assign  RTL__near_mem__WILL_FIRE_server_reset_request_put = RTL__near_mem__EN_server_reset_request_put ; 
  assign  RTL__near_mem__RDY_server_reset_response_get = RTL__near_mem__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__CAN_FIRE_server_reset_response_get = RTL__near_mem__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__WILL_FIRE_server_reset_response_get = RTL__near_mem__EN_server_reset_response_get ; 
  assign  RTL__near_mem__CAN_FIRE_imem_req =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_imem_req = RTL__near_mem__EN_imem_req ; 
  assign  RTL__near_mem__imem_valid = RTL__near_mem__icache$valid ; 
  assign  RTL__near_mem__imem_is_i32_not_i16 =1'd1; 
  assign  RTL__near_mem__imem_pc = RTL__near_mem__icache$addr ; 
  assign  RTL__near_mem__imem_instr ={7'b0,5'bx,5'bx,3'b0,5'bx,7'b0110011}; 
  assign  RTL__near_mem__imem_exc = RTL__near_mem__icache$exc ; 
  assign  RTL__near_mem__imem_exc_code = RTL__near_mem__icache$exc_code ; 
  assign  RTL__near_mem__imem_tval = RTL__near_mem__icache$addr ; 
  assign  RTL__near_mem__imem_master_awvalid = RTL__near_mem__icache$mem_master_awvalid ; 
  assign  RTL__near_mem__imem_master_awid = RTL__near_mem__icache$mem_master_awid ; 
  assign  RTL__near_mem__imem_master_awaddr = RTL__near_mem__icache$mem_master_awaddr ; 
  assign  RTL__near_mem__imem_master_awlen = RTL__near_mem__icache$mem_master_awlen ; 
  assign  RTL__near_mem__imem_master_awsize = RTL__near_mem__icache$mem_master_awsize ; 
  assign  RTL__near_mem__imem_master_awburst = RTL__near_mem__icache$mem_master_awburst ; 
  assign  RTL__near_mem__imem_master_awlock = RTL__near_mem__icache$mem_master_awlock ; 
  assign  RTL__near_mem__imem_master_awcache = RTL__near_mem__icache$mem_master_awcache ; 
  assign  RTL__near_mem__imem_master_awprot = RTL__near_mem__icache$mem_master_awprot ; 
  assign  RTL__near_mem__imem_master_awqos = RTL__near_mem__icache$mem_master_awqos ; 
  assign  RTL__near_mem__imem_master_awregion = RTL__near_mem__icache$mem_master_awregion ; 
  assign  RTL__near_mem__CAN_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL__near_mem__imem_master_wvalid = RTL__near_mem__icache$mem_master_wvalid ; 
  assign  RTL__near_mem__imem_master_wdata = RTL__near_mem__icache$mem_master_wdata ; 
  assign  RTL__near_mem__imem_master_wstrb = RTL__near_mem__icache$mem_master_wstrb ; 
  assign  RTL__near_mem__imem_master_wlast = RTL__near_mem__icache$mem_master_wlast ; 
  assign  RTL__near_mem__CAN_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL__near_mem__CAN_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__imem_master_bready = RTL__near_mem__icache$mem_master_bready ; 
  assign  RTL__near_mem__imem_master_arvalid = RTL__near_mem__icache$mem_master_arvalid ; 
  assign  RTL__near_mem__imem_master_arid = RTL__near_mem__icache$mem_master_arid ; 
  assign  RTL__near_mem__imem_master_araddr = RTL__near_mem__icache$mem_master_araddr ; 
  assign  RTL__near_mem__imem_master_arlen = RTL__near_mem__icache$mem_master_arlen ; 
  assign  RTL__near_mem__imem_master_arsize = RTL__near_mem__icache$mem_master_arsize ; 
  assign  RTL__near_mem__imem_master_arburst = RTL__near_mem__icache$mem_master_arburst ; 
  assign  RTL__near_mem__imem_master_arlock = RTL__near_mem__icache$mem_master_arlock ; 
  assign  RTL__near_mem__imem_master_arcache = RTL__near_mem__icache$mem_master_arcache ; 
  assign  RTL__near_mem__imem_master_arprot = RTL__near_mem__icache$mem_master_arprot ; 
  assign  RTL__near_mem__imem_master_arqos = RTL__near_mem__icache$mem_master_arqos ; 
  assign  RTL__near_mem__imem_master_arregion = RTL__near_mem__icache$mem_master_arregion ; 
  assign  RTL__near_mem__CAN_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL__near_mem__CAN_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__imem_master_rready = RTL__near_mem__icache$mem_master_rready ; 
  assign  RTL__near_mem__CAN_FIRE_dmem_req =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_dmem_req = RTL__near_mem__EN_dmem_req ; 
  assign  RTL__near_mem__dmem_valid = RTL__near_mem__dcache$valid ; 
  assign  RTL__near_mem__dmem_word64 = RTL__near_mem__dcache$word64 ; 
  assign  RTL__near_mem__dmem_st_amo_val =64'hAAAAAAAAAAAAAAAA; 
  assign  RTL__near_mem__dmem_exc = RTL__near_mem__dcache$exc ; 
  assign  RTL__near_mem__dmem_exc_code = RTL__near_mem__dcache$exc_code ; 
  assign  RTL__near_mem__dmem_master_awvalid = RTL__near_mem__dcache$mem_master_awvalid ; 
  assign  RTL__near_mem__dmem_master_awid = RTL__near_mem__dcache$mem_master_awid ; 
  assign  RTL__near_mem__dmem_master_awaddr = RTL__near_mem__dcache$mem_master_awaddr ; 
  assign  RTL__near_mem__dmem_master_awlen = RTL__near_mem__dcache$mem_master_awlen ; 
  assign  RTL__near_mem__dmem_master_awsize = RTL__near_mem__dcache$mem_master_awsize ; 
  assign  RTL__near_mem__dmem_master_awburst = RTL__near_mem__dcache$mem_master_awburst ; 
  assign  RTL__near_mem__dmem_master_awlock = RTL__near_mem__dcache$mem_master_awlock ; 
  assign  RTL__near_mem__dmem_master_awcache = RTL__near_mem__dcache$mem_master_awcache ; 
  assign  RTL__near_mem__dmem_master_awprot = RTL__near_mem__dcache$mem_master_awprot ; 
  assign  RTL__near_mem__dmem_master_awqos = RTL__near_mem__dcache$mem_master_awqos ; 
  assign  RTL__near_mem__dmem_master_awregion = RTL__near_mem__dcache$mem_master_awregion ; 
  assign  RTL__near_mem__CAN_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL__near_mem__dmem_master_wvalid = RTL__near_mem__dcache$mem_master_wvalid ; 
  assign  RTL__near_mem__dmem_master_wdata = RTL__near_mem__dcache$mem_master_wdata ; 
  assign  RTL__near_mem__dmem_master_wstrb = RTL__near_mem__dcache$mem_master_wstrb ; 
  assign  RTL__near_mem__dmem_master_wlast = RTL__near_mem__dcache$mem_master_wlast ; 
  assign  RTL__near_mem__CAN_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL__near_mem__CAN_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__dmem_master_bready = RTL__near_mem__dcache$mem_master_bready ; 
  assign  RTL__near_mem__dmem_master_arvalid = RTL__near_mem__dcache$mem_master_arvalid ; 
  assign  RTL__near_mem__dmem_master_arid = RTL__near_mem__dcache$mem_master_arid ; 
  assign  RTL__near_mem__dmem_master_araddr = RTL__near_mem__dcache$mem_master_araddr ; 
  assign  RTL__near_mem__dmem_master_arlen = RTL__near_mem__dcache$mem_master_arlen ; 
  assign  RTL__near_mem__dmem_master_arsize = RTL__near_mem__dcache$mem_master_arsize ; 
  assign  RTL__near_mem__dmem_master_arburst = RTL__near_mem__dcache$mem_master_arburst ; 
  assign  RTL__near_mem__dmem_master_arlock = RTL__near_mem__dcache$mem_master_arlock ; 
  assign  RTL__near_mem__dmem_master_arcache = RTL__near_mem__dcache$mem_master_arcache ; 
  assign  RTL__near_mem__dmem_master_arprot = RTL__near_mem__dcache$mem_master_arprot ; 
  assign  RTL__near_mem__dmem_master_arqos = RTL__near_mem__dcache$mem_master_arqos ; 
  assign  RTL__near_mem__dmem_master_arregion = RTL__near_mem__dcache$mem_master_arregion ; 
  assign  RTL__near_mem__CAN_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL__near_mem__CAN_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__dmem_master_rready = RTL__near_mem__dcache$mem_master_rready ; 
  assign  RTL__near_mem__RDY_server_fence_i_request_put = RTL__near_mem__dcache$RDY_server_flush_request_put && RTL__near_mem__icache$RDY_server_flush_request_put ; 
  assign  RTL__near_mem__CAN_FIRE_server_fence_i_request_put = RTL__near_mem__dcache$RDY_server_flush_request_put && RTL__near_mem__icache$RDY_server_flush_request_put ; 
  assign  RTL__near_mem__WILL_FIRE_server_fence_i_request_put = RTL__near_mem__EN_server_fence_i_request_put ; 
  assign  RTL__near_mem__RDY_server_fence_i_response_get = RTL__near_mem__dcache$RDY_server_flush_response_get && RTL__near_mem__icache$RDY_server_flush_response_get ; 
  assign  RTL__near_mem__CAN_FIRE_server_fence_i_response_get = RTL__near_mem__dcache$RDY_server_flush_response_get && RTL__near_mem__icache$RDY_server_flush_response_get ; 
  assign  RTL__near_mem__WILL_FIRE_server_fence_i_response_get = RTL__near_mem__EN_server_fence_i_response_get ; 
  assign  RTL__near_mem__RDY_server_fence_request_put = RTL__near_mem__dcache$RDY_server_flush_request_put ; 
  assign  RTL__near_mem__CAN_FIRE_server_fence_request_put = RTL__near_mem__dcache$RDY_server_flush_request_put ; 
  assign  RTL__near_mem__WILL_FIRE_server_fence_request_put = RTL__near_mem__EN_server_fence_request_put ; 
  assign  RTL__near_mem__RDY_server_fence_response_get = RTL__near_mem__dcache$RDY_server_flush_response_get ; 
  assign  RTL__near_mem__CAN_FIRE_server_fence_response_get = RTL__near_mem__dcache$RDY_server_flush_response_get ; 
  assign  RTL__near_mem__WILL_FIRE_server_fence_response_get = RTL__near_mem__EN_server_fence_response_get ; 
  assign  RTL__near_mem__RDY_sfence_vma =1'd1; 
  assign  RTL__near_mem__CAN_FIRE_sfence_vma =1'd1; 
  assign  RTL__near_mem__WILL_FIRE_sfence_vma = RTL__near_mem__EN_sfence_vma ;  
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire[31:0] RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire[31:0] RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL__near_mem__dcache__CLK;
    wire RTL__near_mem__dcache__RST_N;
    wire[3:0] RTL__near_mem__dcache__set_verbosity_verbosity;
    wire RTL__near_mem__dcache__EN_set_verbosity;
    wire RTL__near_mem__dcache__RDY_set_verbosity;
    wire RTL__near_mem__dcache__EN_server_reset_request_put;
    wire RTL__near_mem__dcache__RDY_server_reset_request_put;
    wire RTL__near_mem__dcache__EN_server_reset_response_get;
    wire RTL__near_mem__dcache__RDY_server_reset_response_get;
    wire RTL__near_mem__dcache__req_op;
    wire[2:0] RTL__near_mem__dcache__req_f3;
    wire[31:0] RTL__near_mem__dcache__req_addr;
    wire[63:0] RTL__near_mem__dcache__req_st_value;
    wire[1:0] RTL__near_mem__dcache__req_priv;
    wire RTL__near_mem__dcache__req_sstatus_SUM;
    wire RTL__near_mem__dcache__req_mstatus_MXR;
    wire[31:0] RTL__near_mem__dcache__req_satp;
    wire RTL__near_mem__dcache__EN_req;
    wire RTL__near_mem__dcache__valid;
    wire[31:0] RTL__near_mem__dcache__addr;
    wire[63:0] RTL__near_mem__dcache__word64;
    wire[63:0] RTL__near_mem__dcache__st_amo_val;
    wire RTL__near_mem__dcache__exc;
    wire[3:0] RTL__near_mem__dcache__exc_code;
    wire RTL__near_mem__dcache__EN_server_flush_request_put;
    wire RTL__near_mem__dcache__RDY_server_flush_request_put;
    wire RTL__near_mem__dcache__EN_server_flush_response_get;
    wire RTL__near_mem__dcache__RDY_server_flush_response_get;
    wire RTL__near_mem__dcache__EN_tlb_flush;
    wire RTL__near_mem__dcache__RDY_tlb_flush;
    wire RTL__near_mem__dcache__mem_master_awvalid;
    wire[3:0] RTL__near_mem__dcache__mem_master_awid;
    wire[63:0] RTL__near_mem__dcache__mem_master_awaddr;
    wire[7:0] RTL__near_mem__dcache__mem_master_awlen;
    wire[2:0] RTL__near_mem__dcache__mem_master_awsize;
    wire[1:0] RTL__near_mem__dcache__mem_master_awburst;
    wire RTL__near_mem__dcache__mem_master_awlock;
    wire[3:0] RTL__near_mem__dcache__mem_master_awcache;
    wire[2:0] RTL__near_mem__dcache__mem_master_awprot;
    wire[3:0] RTL__near_mem__dcache__mem_master_awqos;
    wire[3:0] RTL__near_mem__dcache__mem_master_awregion;
    wire RTL__near_mem__dcache__mem_master_awready;
    wire RTL__near_mem__dcache__mem_master_wvalid;
    wire[63:0] RTL__near_mem__dcache__mem_master_wdata;
    wire[7:0] RTL__near_mem__dcache__mem_master_wstrb;
    wire RTL__near_mem__dcache__mem_master_wlast;
    wire RTL__near_mem__dcache__mem_master_wready;
    wire RTL__near_mem__dcache__mem_master_bvalid;
    wire[3:0] RTL__near_mem__dcache__mem_master_bid;
    wire[1:0] RTL__near_mem__dcache__mem_master_bresp;
    wire RTL__near_mem__dcache__mem_master_bready;
    wire RTL__near_mem__dcache__mem_master_arvalid;
    wire[3:0] RTL__near_mem__icache__mem_master_arid;
    wire[63:0] RTL__near_mem__icache__mem_master_araddr;
    wire[7:0] RTL__near_mem__icache__mem_master_arlen;
    wire[2:0] RTL__near_mem__icache__mem_master_arsize;
    wire[1:0] RTL__near_mem__icache__mem_master_arburst;
    wire RTL__near_mem__icache__mem_master_arlock;
    wire[3:0] RTL__near_mem__icache__mem_master_arcache;
    wire[2:0] RTL__near_mem__icache__mem_master_arprot;
    wire[3:0] RTL__near_mem__icache__mem_master_arqos;
    wire[3:0] RTL__near_mem__icache__mem_master_arregion;
    wire RTL__near_mem__icache__mem_master_arready;
    wire RTL__near_mem__icache__mem_master_rvalid;
    wire[3:0] RTL__near_mem__icache__mem_master_rid;
    wire[63:0] RTL__near_mem__icache__mem_master_rdata;
    wire[1:0] RTL__near_mem__icache__mem_master_rresp;
    wire RTL__near_mem__icache__mem_master_rlast;
    wire RTL__near_mem__icache__mem_master_rready;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire[31:0] RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire[31:0] RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL__near_mem__icache__CLK;
    wire RTL__near_mem__icache__RST_N;
    wire[3:0] RTL__near_mem__icache__set_verbosity_verbosity;
    wire RTL__near_mem__icache__EN_set_verbosity;
    wire RTL__near_mem__icache__RDY_set_verbosity;
    wire RTL__near_mem__icache__EN_server_reset_request_put;
    wire RTL__near_mem__icache__RDY_server_reset_request_put;
    wire RTL__near_mem__icache__EN_server_reset_response_get;
    wire RTL__near_mem__icache__RDY_server_reset_response_get;
    wire RTL__near_mem__icache__req_op;
    wire[2:0] RTL__near_mem__icache__req_f3;
    wire[31:0] RTL__near_mem__icache__req_addr;
    wire[63:0] RTL__near_mem__icache__req_st_value;
    wire[1:0] RTL__near_mem__icache__req_priv;
    wire RTL__near_mem__icache__req_sstatus_SUM;
    wire RTL__near_mem__icache__req_mstatus_MXR;
    wire[31:0] RTL__near_mem__icache__req_satp;
    wire RTL__near_mem__icache__EN_req;
    wire RTL__near_mem__icache__valid;
    wire[31:0] RTL__near_mem__icache__addr;
    wire[63:0] RTL__near_mem__icache__word64;
    wire[63:0] RTL__near_mem__icache__st_amo_val;
    wire RTL__near_mem__icache__exc;
    wire[3:0] RTL__near_mem__icache__exc_code;
    wire RTL__near_mem__icache__EN_server_flush_request_put;
    wire RTL__near_mem__icache__RDY_server_flush_request_put;
    wire RTL__near_mem__icache__EN_server_flush_response_get;
    wire RTL__near_mem__icache__RDY_server_flush_response_get;
    wire RTL__near_mem__icache__EN_tlb_flush;
    wire RTL__near_mem__icache__RDY_tlb_flush;
    wire RTL__near_mem__icache__mem_master_awvalid;
    wire[3:0] RTL__near_mem__icache__mem_master_awid;
    wire[63:0] RTL__near_mem__icache__mem_master_awaddr;
    wire[7:0] RTL__near_mem__icache__mem_master_awlen;
    wire[2:0] RTL__near_mem__icache__mem_master_awsize;

    parameter RTL__near_mem__dcache__dmem_not_imem =1'b0; reg[63:0] RTL__near_mem__dcache__word64 ; 
    wire[63:0] RTL__near_mem__dcache__mem_master_araddr , RTL__near_mem__dcache__mem_master_awaddr , RTL__near_mem__dcache__mem_master_wdata , RTL__near_mem__dcache__st_amo_val ; 
    wire[31:0] RTL__near_mem__dcache__addr ; 
    wire[7:0] RTL__near_mem__dcache__mem_master_arlen , RTL__near_mem__dcache__mem_master_awlen , RTL__near_mem__dcache__mem_master_wstrb ; 
    wire[3:0] RTL__near_mem__dcache__exc_code , RTL__near_mem__dcache__mem_master_arcache , RTL__near_mem__dcache__mem_master_arid , RTL__near_mem__dcache__mem_master_arqos , RTL__near_mem__dcache__mem_master_arregion , RTL__near_mem__dcache__mem_master_awcache , RTL__near_mem__dcache__mem_master_awid , RTL__near_mem__dcache__mem_master_awqos , RTL__near_mem__dcache__mem_master_awregion ; 
    wire[2:0] RTL__near_mem__dcache__mem_master_arprot , RTL__near_mem__dcache__mem_master_arsize , RTL__near_mem__dcache__mem_master_awprot , RTL__near_mem__dcache__mem_master_awsize ; 
    wire[1:0] RTL__near_mem__dcache__mem_master_arburst , RTL__near_mem__dcache__mem_master_awburst ; 
    wire RTL__near_mem__dcache__RDY_server_flush_request_put , RTL__near_mem__dcache__RDY_server_flush_response_get , RTL__near_mem__dcache__RDY_server_reset_request_put , RTL__near_mem__dcache__RDY_server_reset_response_get , RTL__near_mem__dcache__RDY_set_verbosity , RTL__near_mem__dcache__RDY_tlb_flush , RTL__near_mem__dcache__exc , RTL__near_mem__dcache__mem_master_arlock , RTL__near_mem__dcache__mem_master_arvalid , RTL__near_mem__dcache__mem_master_awlock , RTL__near_mem__dcache__mem_master_awvalid , RTL__near_mem__dcache__mem_master_bready , RTL__near_mem__dcache__mem_master_rready , RTL__near_mem__dcache__mem_master_wlast , RTL__near_mem__dcache__mem_master_wvalid , RTL__near_mem__dcache__valid ; 
    wire[3:0] RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port0__write_1 , RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port1__write_1 , RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port2__read , RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port3__read ; 
    wire RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$EN_port2__write , RTL__near_mem__dcache__dw_valid$whas ; reg[3:0] RTL__near_mem__dcache__cfg_verbosity ; 
    wire[3:0] RTL__near_mem__dcache__cfg_verbosity$D_IN ; 
    wire RTL__near_mem__dcache__cfg_verbosity$EN ; reg[3:0] RTL__near_mem__dcache__ctr_wr_rsps_pending_crg ; 
    wire[3:0] RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$D_IN ; 
    wire RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$EN ; reg[31:0] RTL__near_mem__dcache__rg_addr ; 
    wire[31:0] RTL__near_mem__dcache__rg_addr$D_IN ; 
    wire RTL__near_mem__dcache__rg_addr$EN ; reg[6:0] RTL__near_mem__dcache__rg_cset_in_cache ; 
    wire[6:0] RTL__near_mem__dcache__rg_cset_in_cache$D_IN ; 
    wire RTL__near_mem__dcache__rg_cset_in_cache$EN ; 
    reg RTL__near_mem__dcache__rg_error_during_refill ; 
    wire RTL__near_mem__dcache__rg_error_during_refill$D_IN , RTL__near_mem__dcache__rg_error_during_refill$EN ; reg[3:0] RTL__near_mem__dcache__rg_exc_code ; reg[3:0] RTL__near_mem__dcache__rg_exc_code$D_IN ; 
    wire RTL__near_mem__dcache__rg_exc_code$EN ; reg[2:0] RTL__near_mem__dcache__rg_f3 ; 
    wire[2:0] RTL__near_mem__dcache__rg_f3$D_IN ; 
    wire RTL__near_mem__dcache__rg_f3$EN ; reg[63:0] RTL__near_mem__dcache__rg_ld_val ; 
    wire[63:0] RTL__near_mem__dcache__rg_ld_val$D_IN ; 
    wire RTL__near_mem__dcache__rg_ld_val$EN ; reg[31:0] RTL__near_mem__dcache__rg_lower_word32 ; 
    wire[31:0] RTL__near_mem__dcache__rg_lower_word32$D_IN ; 
    wire RTL__near_mem__dcache__rg_lower_word32$EN ; 
    reg RTL__near_mem__dcache__rg_lower_word32_full ; 
    wire RTL__near_mem__dcache__rg_lower_word32_full$D_IN , RTL__near_mem__dcache__rg_lower_word32_full$EN ; 
    reg RTL__near_mem__dcache__rg_op ; 
    wire RTL__near_mem__dcache__rg_op$D_IN , RTL__near_mem__dcache__rg_op$EN ; reg[31:0] RTL__near_mem__dcache__rg_pa ; 
    wire[31:0] RTL__near_mem__dcache__rg_pa$D_IN ; 
    wire RTL__near_mem__dcache__rg_pa$EN ; reg[31:0] RTL__near_mem__dcache__rg_pte_pa ; 
    wire[31:0] RTL__near_mem__dcache__rg_pte_pa$D_IN ; 
    wire RTL__near_mem__dcache__rg_pte_pa$EN ; reg[63:0] RTL__near_mem__dcache__rg_st_amo_val ; 
    wire[63:0] RTL__near_mem__dcache__rg_st_amo_val$D_IN ; 
    wire RTL__near_mem__dcache__rg_st_amo_val$EN ; reg[3:0] RTL__near_mem__dcache__rg_state ; reg[3:0] RTL__near_mem__dcache__rg_state$D_IN ; 
    wire RTL__near_mem__dcache__rg_state$EN ; reg[8:0] RTL__near_mem__dcache__rg_word64_set_in_cache ; 
    wire[8:0] RTL__near_mem__dcache__rg_word64_set_in_cache$D_IN ; 
    wire RTL__near_mem__dcache__rg_word64_set_in_cache$EN ; 
    wire[98:0] RTL__near_mem__dcache__f_fabric_write_reqs$D_IN , RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT ; 
    wire RTL__near_mem__dcache__f_fabric_write_reqs$CLR , RTL__near_mem__dcache__f_fabric_write_reqs$DEQ , RTL__near_mem__dcache__f_fabric_write_reqs$EMPTY_N , RTL__near_mem__dcache__f_fabric_write_reqs$ENQ , RTL__near_mem__dcache__f_fabric_write_reqs$FULL_N ; 
    wire RTL__near_mem__dcache__f_reset_reqs$CLR , RTL__near_mem__dcache__f_reset_reqs$DEQ , RTL__near_mem__dcache__f_reset_reqs$D_IN , RTL__near_mem__dcache__f_reset_reqs$D_OUT , RTL__near_mem__dcache__f_reset_reqs$EMPTY_N , RTL__near_mem__dcache__f_reset_reqs$ENQ , RTL__near_mem__dcache__f_reset_reqs$FULL_N ; 
    wire RTL__near_mem__dcache__f_reset_rsps$CLR , RTL__near_mem__dcache__f_reset_rsps$DEQ , RTL__near_mem__dcache__f_reset_rsps$D_IN , RTL__near_mem__dcache__f_reset_rsps$D_OUT , RTL__near_mem__dcache__f_reset_rsps$EMPTY_N , RTL__near_mem__dcache__f_reset_rsps$ENQ , RTL__near_mem__dcache__f_reset_rsps$FULL_N ; 
    wire[96:0] RTL__near_mem__dcache__master_xactor_f_rd_addr$D_IN , RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT ; 
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr$CLR , RTL__near_mem__dcache__master_xactor_f_rd_addr$DEQ , RTL__near_mem__dcache__master_xactor_f_rd_addr$EMPTY_N , RTL__near_mem__dcache__master_xactor_f_rd_addr$ENQ , RTL__near_mem__dcache__master_xactor_f_rd_addr$FULL_N ; 
    wire[70:0] RTL__near_mem__dcache__master_xactor_f_rd_data$D_IN , RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT ; 
    wire RTL__near_mem__dcache__master_xactor_f_rd_data$CLR , RTL__near_mem__dcache__master_xactor_f_rd_data$DEQ , RTL__near_mem__dcache__master_xactor_f_rd_data$EMPTY_N , RTL__near_mem__dcache__master_xactor_f_rd_data$ENQ , RTL__near_mem__dcache__master_xactor_f_rd_data$FULL_N ; 
    wire[96:0] RTL__near_mem__dcache__master_xactor_f_wr_addr$D_IN , RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr$CLR , RTL__near_mem__dcache__master_xactor_f_wr_addr$DEQ , RTL__near_mem__dcache__master_xactor_f_wr_addr$EMPTY_N , RTL__near_mem__dcache__master_xactor_f_wr_addr$ENQ , RTL__near_mem__dcache__master_xactor_f_wr_addr$FULL_N ; 
    wire[72:0] RTL__near_mem__dcache__master_xactor_f_wr_data$D_IN , RTL__near_mem__dcache__master_xactor_f_wr_data$D_OUT ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_data$CLR , RTL__near_mem__dcache__master_xactor_f_wr_data$DEQ , RTL__near_mem__dcache__master_xactor_f_wr_data$EMPTY_N , RTL__near_mem__dcache__master_xactor_f_wr_data$ENQ , RTL__near_mem__dcache__master_xactor_f_wr_data$FULL_N ; 
    wire[5:0] RTL__near_mem__dcache__master_xactor_f_wr_resp$D_IN , RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp$CLR , RTL__near_mem__dcache__master_xactor_f_wr_resp$DEQ , RTL__near_mem__dcache__master_xactor_f_wr_resp$EMPTY_N , RTL__near_mem__dcache__master_xactor_f_wr_resp$ENQ , RTL__near_mem__dcache__master_xactor_f_wr_resp$FULL_N ; 
    wire[22:0] RTL__near_mem__dcache__ram_state_and_ctag_cset$DIA , RTL__near_mem__dcache__ram_state_and_ctag_cset$DIB , RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB ; 
    wire[6:0] RTL__near_mem__dcache__ram_state_and_ctag_cset$ADDRA , RTL__near_mem__dcache__ram_state_and_ctag_cset$ADDRB ; 
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset$ENA , RTL__near_mem__dcache__ram_state_and_ctag_cset$ENB , RTL__near_mem__dcache__ram_state_and_ctag_cset$WEA , RTL__near_mem__dcache__ram_state_and_ctag_cset$WEB ; reg[63:0] RTL__near_mem__dcache__ram_word64_set$DIB ; reg[8:0] RTL__near_mem__dcache__ram_word64_set$ADDRB ; 
    wire[63:0] RTL__near_mem__dcache__ram_word64_set$DIA , RTL__near_mem__dcache__ram_word64_set$DOB ; 
    wire[8:0] RTL__near_mem__dcache__ram_word64_set$ADDRA ; 
    wire RTL__near_mem__dcache__ram_word64_set$ENA , RTL__near_mem__dcache__ram_word64_set$ENB , RTL__near_mem__dcache__ram_word64_set$WEA , RTL__near_mem__dcache__ram_word64_set$WEB ; 
    wire[63:0] RTL__near_mem__dcache__soc_map$m_is_IO_addr_addr , RTL__near_mem__dcache__soc_map$m_is_mem_addr_addr , RTL__near_mem__dcache__soc_map$m_is_near_mem_IO_addr_addr ; 
    wire RTL__near_mem__dcache__soc_map$m_is_mem_addr ; 
    wire RTL__near_mem__dcache__CAN_FIRE_RL_rl_ST_AMO_response , RTL__near_mem__dcache__CAN_FIRE_RL_rl_cache_refill_rsps_loop , RTL__near_mem__dcache__CAN_FIRE_RL_rl_discard_write_rsp , RTL__near_mem__dcache__CAN_FIRE_RL_rl_drive_exception_rsp , RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req , RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_read_req , RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_read_rsp , RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_write_req , RTL__near_mem__dcache__CAN_FIRE_RL_rl_maintain_io_read_rsp , RTL__near_mem__dcache__CAN_FIRE_RL_rl_probe_and_immed_rsp , RTL__near_mem__dcache__CAN_FIRE_RL_rl_rereq , RTL__near_mem__dcache__CAN_FIRE_RL_rl_reset , RTL__near_mem__dcache__CAN_FIRE_RL_rl_start_cache_refill , RTL__near_mem__dcache__CAN_FIRE_RL_rl_start_reset , RTL__near_mem__dcache__CAN_FIRE_mem_master_m_arready , RTL__near_mem__dcache__CAN_FIRE_mem_master_m_awready , RTL__near_mem__dcache__CAN_FIRE_mem_master_m_bvalid , RTL__near_mem__dcache__CAN_FIRE_mem_master_m_rvalid , RTL__near_mem__dcache__CAN_FIRE_mem_master_m_wready , RTL__near_mem__dcache__CAN_FIRE_req , RTL__near_mem__dcache__CAN_FIRE_server_flush_request_put , RTL__near_mem__dcache__CAN_FIRE_server_flush_response_get , RTL__near_mem__dcache__CAN_FIRE_server_reset_request_put , RTL__near_mem__dcache__CAN_FIRE_server_reset_response_get , RTL__near_mem__dcache__CAN_FIRE_set_verbosity , RTL__near_mem__dcache__CAN_FIRE_tlb_flush , RTL__near_mem__dcache__WILL_FIRE_RL_rl_ST_AMO_response , RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop , RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp , RTL__near_mem__dcache__WILL_FIRE_RL_rl_drive_exception_rsp , RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req , RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req , RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp , RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req , RTL__near_mem__dcache__WILL_FIRE_RL_rl_maintain_io_read_rsp , RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp , RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq , RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset , RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill , RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset , RTL__near_mem__dcache__WILL_FIRE_mem_master_m_arready , RTL__near_mem__dcache__WILL_FIRE_mem_master_m_awready , RTL__near_mem__dcache__WILL_FIRE_mem_master_m_bvalid , RTL__near_mem__dcache__WILL_FIRE_mem_master_m_rvalid , RTL__near_mem__dcache__WILL_FIRE_mem_master_m_wready , RTL__near_mem__dcache__WILL_FIRE_req , RTL__near_mem__dcache__WILL_FIRE_server_flush_request_put , RTL__near_mem__dcache__WILL_FIRE_server_flush_response_get , RTL__near_mem__dcache__WILL_FIRE_server_reset_request_put , RTL__near_mem__dcache__WILL_FIRE_server_reset_response_get , RTL__near_mem__dcache__WILL_FIRE_set_verbosity , RTL__near_mem__dcache__WILL_FIRE_tlb_flush ; reg[63:0] RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2 ; 
    wire[98:0] RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__VAL_1 , RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
    wire[96:0] RTL__near_mem__dcache__MUX_master_xactor_f_rd_addr$enq_1__VAL_1 , RTL__near_mem__dcache__MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
    wire[22:0] RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ; 
    wire[8:0] RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_2 , RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_4 ; 
    wire[6:0] RTL__near_mem__dcache__MUX_rg_cset_in_cache$write_1__VAL_1 ; 
    wire[3:0] RTL__near_mem__dcache__MUX_rg_exc_code$write_1__VAL_1 , RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_1 , RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_4 , RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_7 , RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_9 ; 
    wire RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_1 , RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_2 , RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_3 , RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__SEL_1 , RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 , RTL__near_mem__dcache__MUX_ram_word64_set$a_put_1__SEL_1 , RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2 , RTL__near_mem__dcache__MUX_rg_error_during_refill$write_1__SEL_1 , RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_1 , RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_2 , RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_10 , RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_2 , RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_3 , RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_7 , RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_9 ; reg[31:0] RTL__near_mem__dcache__v__h2948 ; reg[31:0] RTL__near_mem__dcache__v__h3848 ; reg[31:0] RTL__near_mem__dcache__v__h3949 ; reg[31:0] RTL__near_mem__dcache__v__h4098 ; reg[31:0] RTL__near_mem__dcache__v__h12540 ; reg[31:0] RTL__near_mem__dcache__v__h14531 ; reg[31:0] RTL__near_mem__dcache__v__h15336 ; reg[31:0] RTL__near_mem__dcache__v__h15578 ; reg[31:0] RTL__near_mem__dcache__v__h17191 ; reg[31:0] RTL__near_mem__dcache__v__h17485 ; reg[31:0] RTL__near_mem__dcache__v__h18585 ; reg[31:0] RTL__near_mem__dcache__v__h18692 ; reg[31:0] RTL__near_mem__dcache__v__h18797 ; reg[31:0] RTL__near_mem__dcache__v__h18877 ; reg[31:0] RTL__near_mem__dcache__v__h19505 ; reg[31:0] RTL__near_mem__dcache__v__h19466 ; reg[31:0] RTL__near_mem__dcache__v__h3483 ; reg[31:0] RTL__near_mem__dcache__v__h19852 ; reg[31:0] RTL__near_mem__dcache__v__h2942 ; reg[31:0] RTL__near_mem__dcache__v__h3477 ; reg[31:0] RTL__near_mem__dcache__v__h3842 ; reg[31:0] RTL__near_mem__dcache__v__h3943 ; reg[31:0] RTL__near_mem__dcache__v__h4092 ; reg[31:0] RTL__near_mem__dcache__v__h12534 ; reg[31:0] RTL__near_mem__dcache__v__h14525 ; reg[31:0] RTL__near_mem__dcache__v__h15330 ; reg[31:0] RTL__near_mem__dcache__v__h15572 ; reg[31:0] RTL__near_mem__dcache__v__h17185 ; reg[31:0] RTL__near_mem__dcache__v__h17479 ; reg[31:0] RTL__near_mem__dcache__v__h18579 ; reg[31:0] RTL__near_mem__dcache__v__h18686 ; reg[31:0] RTL__near_mem__dcache__v__h18791 ; reg[31:0] RTL__near_mem__dcache__v__h18871 ; reg[31:0] RTL__near_mem__dcache__v__h19460 ; reg[31:0] RTL__near_mem__dcache__v__h19499 ; reg[31:0] RTL__near_mem__dcache__v__h19846 ; reg[63:0] RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 , RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 , RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 , RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 , RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 , RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 , RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 , RTL__near_mem__dcache__ld_val__h17594 , RTL__near_mem__dcache__mem_req_wr_data_wdata__h2699 ; reg[7:0] RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700 ; reg[2:0] RTL__near_mem__dcache__value__h17372 , RTL__near_mem__dcache__x__h2520 ; 
    wire[63:0] RTL__near_mem__dcache___theResult___snd_fst__h2707 , RTL__near_mem__dcache__cline_fabric_addr__h14584 , RTL__near_mem__dcache__fabric_addr__h17243 , RTL__near_mem__dcache__mem_req_wr_addr_awaddr__h2473 , RTL__near_mem__dcache__result__h11657 , RTL__near_mem__dcache__result__h11685 , RTL__near_mem__dcache__result__h11713 , RTL__near_mem__dcache__result__h11741 , RTL__near_mem__dcache__result__h11769 , RTL__near_mem__dcache__result__h11797 , RTL__near_mem__dcache__result__h11825 , RTL__near_mem__dcache__result__h11870 , RTL__near_mem__dcache__result__h11898 , RTL__near_mem__dcache__result__h11926 , RTL__near_mem__dcache__result__h11954 , RTL__near_mem__dcache__result__h11982 , RTL__near_mem__dcache__result__h12010 , RTL__near_mem__dcache__result__h12038 , RTL__near_mem__dcache__result__h12066 , RTL__near_mem__dcache__result__h12111 , RTL__near_mem__dcache__result__h12139 , RTL__near_mem__dcache__result__h12167 , RTL__near_mem__dcache__result__h12195 , RTL__near_mem__dcache__result__h12236 , RTL__near_mem__dcache__result__h12264 , RTL__near_mem__dcache__result__h12292 , RTL__near_mem__dcache__result__h12320 , RTL__near_mem__dcache__result__h12361 , RTL__near_mem__dcache__result__h12389 , RTL__near_mem__dcache__result__h12428 , RTL__near_mem__dcache__result__h12456 , RTL__near_mem__dcache__result__h17654 , RTL__near_mem__dcache__result__h17684 , RTL__near_mem__dcache__result__h17711 , RTL__near_mem__dcache__result__h17738 , RTL__near_mem__dcache__result__h17765 , RTL__near_mem__dcache__result__h17792 , RTL__near_mem__dcache__result__h17819 , RTL__near_mem__dcache__result__h17846 , RTL__near_mem__dcache__result__h17890 , RTL__near_mem__dcache__result__h17917 , RTL__near_mem__dcache__result__h17944 , RTL__near_mem__dcache__result__h17971 , RTL__near_mem__dcache__result__h17998 , RTL__near_mem__dcache__result__h18025 , RTL__near_mem__dcache__result__h18052 , RTL__near_mem__dcache__result__h18079 , RTL__near_mem__dcache__result__h18123 , RTL__near_mem__dcache__result__h18150 , RTL__near_mem__dcache__result__h18177 , RTL__near_mem__dcache__result__h18204 , RTL__near_mem__dcache__result__h18244 , RTL__near_mem__dcache__result__h18271 , RTL__near_mem__dcache__result__h18298 , RTL__near_mem__dcache__result__h18325 , RTL__near_mem__dcache__result__h18365 , RTL__near_mem__dcache__result__h18392 , RTL__near_mem__dcache__result__h18430 , RTL__near_mem__dcache__result__h18457 , RTL__near_mem__dcache__result__h5301 , RTL__near_mem__dcache__word64__h5094 , RTL__near_mem__dcache__y__h5337 ; 
    wire[31:0] RTL__near_mem__dcache__cline_addr__h14583 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 , RTL__near_mem__dcache__word64094_BITS_31_TO_0__q17 , RTL__near_mem__dcache__word64094_BITS_63_TO_32__q24 ; 
    wire[21:0] RTL__near_mem__dcache__pa_ctag__h4952 ; 
    wire[15:0] RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 , RTL__near_mem__dcache__word64094_BITS_15_TO_0__q16 , RTL__near_mem__dcache__word64094_BITS_31_TO_16__q20 , RTL__near_mem__dcache__word64094_BITS_47_TO_32__q23 , RTL__near_mem__dcache__word64094_BITS_63_TO_48__q27 ; 
    wire[7:0] RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 , RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 , RTL__near_mem__dcache__strobe64__h2637 , RTL__near_mem__dcache__strobe64__h2639 , RTL__near_mem__dcache__strobe64__h2641 , RTL__near_mem__dcache__word64094_BITS_15_TO_8__q18 , RTL__near_mem__dcache__word64094_BITS_23_TO_16__q19 , RTL__near_mem__dcache__word64094_BITS_31_TO_24__q21 , RTL__near_mem__dcache__word64094_BITS_39_TO_32__q22 , RTL__near_mem__dcache__word64094_BITS_47_TO_40__q25 , RTL__near_mem__dcache__word64094_BITS_55_TO_48__q26 , RTL__near_mem__dcache__word64094_BITS_63_TO_56__q28 , RTL__near_mem__dcache__word64094_BITS_7_TO_0__q15 ; 
    wire[5:0] RTL__near_mem__dcache__shift_bits__h2487 ; 
    wire[3:0] RTL__near_mem__dcache__access_exc_code__h2256 , RTL__near_mem__dcache__b__h14485 ; 
    wire RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 , RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 , RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 , RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 , RTL__near_mem__dcache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 , RTL__near_mem__dcache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 , RTL__near_mem__dcache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 , RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 , RTL__near_mem__dcache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 , RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 ; 
  assign  RTL__near_mem__dcache__RDY_set_verbosity =1'd1; 
  assign  RTL__near_mem__dcache__CAN_FIRE_set_verbosity =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_set_verbosity = RTL__near_mem__dcache__EN_set_verbosity ; 
  assign  RTL__near_mem__dcache__RDY_server_reset_request_put = RTL__near_mem__dcache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_server_reset_request_put = RTL__near_mem__dcache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_server_reset_request_put = RTL__near_mem__dcache__EN_server_reset_request_put ; 
  assign  RTL__near_mem__dcache__RDY_server_reset_response_get =! RTL__near_mem__dcache__f_reset_rsps$D_OUT && RTL__near_mem__dcache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_server_reset_response_get =! RTL__near_mem__dcache__f_reset_rsps$D_OUT && RTL__near_mem__dcache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_server_reset_response_get = RTL__near_mem__dcache__EN_server_reset_response_get ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_req =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_req = RTL__near_mem__dcache__EN_req ; 
  assign  RTL__near_mem__dcache__valid = RTL__near_mem__dcache__dw_valid$whas ; 
  assign  RTL__near_mem__dcache__addr = RTL__near_mem__dcache__rg_addr ; 
  always @(       RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_1                    or   RTL__near_mem__dcache__ld_val__h17594              or   RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_2             or   RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2            or   RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_3           or   RTL__near_mem__dcache__rg_ld_val  )
         begin 
             case (1'b1) 
              RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_1  : 
                  RTL__near_mem__dcache__word64  = RTL__near_mem__dcache__ld_val__h17594 ; 
              RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_2  : 
                  RTL__near_mem__dcache__word64  = RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2 ; 
              RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_3  : 
                  RTL__near_mem__dcache__word64  = RTL__near_mem__dcache__rg_ld_val ;
              default : 
                  RTL__near_mem__dcache__word64  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL__near_mem__dcache__st_amo_val = RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_2  ? 64'd0: RTL__near_mem__dcache__rg_st_amo_val ; 
  assign  RTL__near_mem__dcache__exc = RTL__near_mem__dcache__rg_state ==4'd4; 
  assign  RTL__near_mem__dcache__exc_code = RTL__near_mem__dcache__rg_exc_code ; 
  assign  RTL__near_mem__dcache__RDY_server_flush_request_put = RTL__near_mem__dcache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_server_flush_request_put = RTL__near_mem__dcache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_server_flush_request_put = RTL__near_mem__dcache__EN_server_flush_request_put ; 
  assign  RTL__near_mem__dcache__RDY_server_flush_response_get = RTL__near_mem__dcache__f_reset_rsps$D_OUT && RTL__near_mem__dcache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_server_flush_response_get = RTL__near_mem__dcache__f_reset_rsps$D_OUT && RTL__near_mem__dcache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_server_flush_response_get = RTL__near_mem__dcache__EN_server_flush_response_get ; 
  assign  RTL__near_mem__dcache__RDY_tlb_flush =1'd1; 
  assign  RTL__near_mem__dcache__CAN_FIRE_tlb_flush =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_tlb_flush = RTL__near_mem__dcache__EN_tlb_flush ; 
  assign  RTL__near_mem__dcache__mem_master_awvalid = RTL__near_mem__dcache__master_xactor_f_wr_addr$EMPTY_N ; 
  assign  RTL__near_mem__dcache__mem_master_awid = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [96:93]; 
  assign  RTL__near_mem__dcache__mem_master_awaddr = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [92:29]; 
  assign  RTL__near_mem__dcache__mem_master_awlen = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [28:21]; 
  assign  RTL__near_mem__dcache__mem_master_awsize = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [20:18]; 
  assign  RTL__near_mem__dcache__mem_master_awburst = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [17:16]; 
  assign  RTL__near_mem__dcache__mem_master_awlock = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [15]; 
  assign  RTL__near_mem__dcache__mem_master_awcache = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [14:11]; 
  assign  RTL__near_mem__dcache__mem_master_awprot = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [10:8]; 
  assign  RTL__near_mem__dcache__mem_master_awqos = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [7:4]; 
  assign  RTL__near_mem__dcache__mem_master_awregion = RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT [3:0]; 
  assign  RTL__near_mem__dcache__CAN_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL__near_mem__dcache__mem_master_wvalid = RTL__near_mem__dcache__master_xactor_f_wr_data$EMPTY_N ; 
  assign  RTL__near_mem__dcache__mem_master_wdata = RTL__near_mem__dcache__master_xactor_f_wr_data$D_OUT [72:9]; 
  assign  RTL__near_mem__dcache__mem_master_wstrb = RTL__near_mem__dcache__master_xactor_f_wr_data$D_OUT [8:1]; 
  assign  RTL__near_mem__dcache__mem_master_wlast = RTL__near_mem__dcache__master_xactor_f_wr_data$D_OUT [0]; 
  assign  RTL__near_mem__dcache__CAN_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL__near_mem__dcache__CAN_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__dcache__mem_master_bready = RTL__near_mem__dcache__master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL__near_mem__dcache__mem_master_arvalid = RTL__near_mem__dcache__master_xactor_f_rd_addr$EMPTY_N ; 
  assign  RTL__near_mem__dcache__mem_master_arid = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [96:93]; 
  assign  RTL__near_mem__dcache__mem_master_araddr = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [92:29]; 
  assign  RTL__near_mem__dcache__mem_master_arlen = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [28:21]; 
  assign  RTL__near_mem__dcache__mem_master_arsize = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [20:18]; 
  assign  RTL__near_mem__dcache__mem_master_arburst = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [17:16]; 
  assign  RTL__near_mem__dcache__mem_master_arlock = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [15]; 
  assign  RTL__near_mem__dcache__mem_master_arcache = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [14:11]; 
  assign  RTL__near_mem__dcache__mem_master_arprot = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [10:8]; 
  assign  RTL__near_mem__dcache__mem_master_arqos = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [7:4]; 
  assign  RTL__near_mem__dcache__mem_master_arregion = RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT [3:0]; 
  assign  RTL__near_mem__dcache__CAN_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL__near_mem__dcache__CAN_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__dcache__mem_master_rready = RTL__near_mem__dcache__master_xactor_f_rd_data$FULL_N ;  
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__f_reset_rsps__CLK;
    wire RTL__near_mem__dcache__f_reset_rsps__RST;
    wire[RTL__near_mem__dcache__f_fabric_write_reqs__width-1:0] RTL__near_mem__dcache__f_reset_rsps__D_IN;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__CLR;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__FULL_N;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__EMPTY_N;
    wire[RTL__near_mem__dcache__f_fabric_write_reqs__width-1:0] RTL__near_mem__dcache__master_xactor_f_rd_addr__D_OUT;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__CLK;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__RST;
    wire[RTL__near_mem__dcache__f_reset_reqs__width-1:0] RTL__near_mem__dcache__master_xactor_f_wr_data__D_IN;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__CLR;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__FULL_N;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__EMPTY_N;
    wire[RTL__near_mem__dcache__f_reset_reqs__width-1:0] RTL__near_mem__dcache__master_xactor_f_wr_data__D_OUT;
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_reqs__CLK;
    wire RTL__near_mem__icache__f_reset_reqs__RST;
    wire[RTL__near_mem__dcache__f_reset_rsps__width-1:0] RTL__near_mem__icache__f_reset_reqs__D_IN;
    wire RTL__near_mem__icache__f_reset_reqs__ENQ;
    wire RTL__near_mem__icache__f_reset_rsps__DEQ;
    wire RTL__near_mem__icache__f_reset_rsps__CLR;
    wire RTL__near_mem__icache__f_reset_rsps__FULL_N;
    wire RTL__near_mem__icache__f_reset_rsps__EMPTY_N;
    wire[RTL__near_mem__dcache__f_reset_rsps__width-1:0] RTL__near_mem__icache__f_reset_rsps__D_OUT;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__CLK;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__RST;
    wire[RTL__near_mem__dcache__master_xactor_f_rd_addr__width-1:0] RTL__near_mem__icache__master_xactor_f_wr_addr__D_IN;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__CLR;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__FULL_N;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__EMPTY_N;
    wire[RTL__near_mem__dcache__master_xactor_f_rd_addr__width-1:0] RTL__near_mem__icache__master_xactor_f_wr_addr__D_OUT;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;

    parameter RTL__near_mem__dcache__f_fabric_write_reqs__width =1; parameter RTL__near_mem__dcache__f_fabric_write_reqs__guarded =1; 
    reg RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
    reg RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; reg[ RTL__near_mem__dcache__f_fabric_write_reqs__width -1:0] RTL__near_mem__dcache__f_fabric_write_reqs__data0_reg ; reg[ RTL__near_mem__dcache__f_fabric_write_reqs__width -1:0] RTL__near_mem__dcache__f_fabric_write_reqs__data1_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__FULL_N = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__EMPTY_N = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__D_OUT = RTL__near_mem__dcache__f_fabric_write_reqs__data0_reg ; 
    wire RTL__near_mem__dcache__f_fabric_write_reqs__d0di =( RTL__near_mem__dcache__f_fabric_write_reqs__ENQ &&! RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg )||( RTL__near_mem__dcache__f_fabric_write_reqs__ENQ && RTL__near_mem__dcache__f_fabric_write_reqs__DEQ && RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ); 
    wire RTL__near_mem__dcache__f_fabric_write_reqs__d0d1 = RTL__near_mem__dcache__f_fabric_write_reqs__DEQ &&! RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
    wire RTL__near_mem__dcache__f_fabric_write_reqs__d0h =((! RTL__near_mem__dcache__f_fabric_write_reqs__DEQ )&&(! RTL__near_mem__dcache__f_fabric_write_reqs__ENQ ))||(! RTL__near_mem__dcache__f_fabric_write_reqs__DEQ && RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg )||(! RTL__near_mem__dcache__f_fabric_write_reqs__ENQ && RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ); 
    wire RTL__near_mem__dcache__f_fabric_write_reqs__d1di = RTL__near_mem__dcache__f_fabric_write_reqs__ENQ & RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__f_fabric_write_reqs__CLK )
         begin 
             if ( RTL__near_mem__dcache__f_fabric_write_reqs__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__f_fabric_write_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__f_fabric_write_reqs__CLR )
                         begin  
                             RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__f_fabric_write_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__f_fabric_write_reqs__ENQ &&! RTL__near_mem__dcache__f_fabric_write_reqs__DEQ )
                             begin  
                                 RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__f_fabric_write_reqs__full_reg  <=! RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__f_fabric_write_reqs__DEQ &&! RTL__near_mem__dcache__f_fabric_write_reqs__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__f_fabric_write_reqs__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg  <=! RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__f_fabric_write_reqs__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__f_fabric_write_reqs__data0_reg  <={ RTL__near_mem__dcache__f_fabric_write_reqs__width { RTL__near_mem__dcache__f_fabric_write_reqs__d0di }}& RTL__near_mem__dcache__f_fabric_write_reqs__D_IN |{ RTL__near_mem__dcache__f_fabric_write_reqs__width { RTL__near_mem__dcache__f_fabric_write_reqs__d0d1 }}& RTL__near_mem__dcache__f_fabric_write_reqs__data1_reg |{ RTL__near_mem__dcache__f_fabric_write_reqs__width { RTL__near_mem__dcache__f_fabric_write_reqs__d0h }}& RTL__near_mem__dcache__f_fabric_write_reqs__data0_reg ; 
                 RTL__near_mem__dcache__f_fabric_write_reqs__data1_reg  <= RTL__near_mem__dcache__f_fabric_write_reqs__d1di  ?  RTL__near_mem__dcache__f_fabric_write_reqs__D_IN : RTL__near_mem__dcache__f_fabric_write_reqs__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__f_fabric_write_reqs__CLK )
         begin : RTL__near_mem__dcache__f_fabric_write_reqs__error_checks 
           reg RTL__near_mem__dcache__f_fabric_write_reqs__deqerror , RTL__near_mem__dcache__f_fabric_write_reqs__enqerror ; 
             RTL__near_mem__dcache__f_fabric_write_reqs__deqerror  =0; 
             RTL__near_mem__dcache__f_fabric_write_reqs__enqerror  =0;
             if ( RTL__near_mem__dcache__f_fabric_write_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg && RTL__near_mem__dcache__f_fabric_write_reqs__DEQ )
                         begin  
                             RTL__near_mem__dcache__f_fabric_write_reqs__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__f_fabric_write_reqs__full_reg && RTL__near_mem__dcache__f_fabric_write_reqs__ENQ &&(! RTL__near_mem__dcache__f_fabric_write_reqs__DEQ || RTL__near_mem__dcache__f_fabric_write_reqs__guarded ))
                         begin  
                             RTL__near_mem__dcache__f_fabric_write_reqs__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__empty_reg ;
    parameter RTL__near_mem__dcache__f_reset_reqs__width =1; parameter RTL__near_mem__dcache__f_reset_reqs__guarded =1; 
    reg RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
    reg RTL__near_mem__dcache__f_reset_reqs__empty_reg ; reg[ RTL__near_mem__dcache__f_reset_reqs__width -1:0] RTL__near_mem__dcache__f_reset_reqs__data0_reg ; reg[ RTL__near_mem__dcache__f_reset_reqs__width -1:0] RTL__near_mem__dcache__f_reset_reqs__data1_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__FULL_N = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__EMPTY_N = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__D_OUT = RTL__near_mem__dcache__f_reset_reqs__data0_reg ; 
    wire RTL__near_mem__dcache__f_reset_reqs__d0di =( RTL__near_mem__dcache__f_reset_reqs__ENQ &&! RTL__near_mem__dcache__f_reset_reqs__empty_reg )||( RTL__near_mem__dcache__f_reset_reqs__ENQ && RTL__near_mem__dcache__f_reset_reqs__DEQ && RTL__near_mem__dcache__f_reset_reqs__full_reg ); 
    wire RTL__near_mem__dcache__f_reset_reqs__d0d1 = RTL__near_mem__dcache__f_reset_reqs__DEQ &&! RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
    wire RTL__near_mem__dcache__f_reset_reqs__d0h =((! RTL__near_mem__dcache__f_reset_reqs__DEQ )&&(! RTL__near_mem__dcache__f_reset_reqs__ENQ ))||(! RTL__near_mem__dcache__f_reset_reqs__DEQ && RTL__near_mem__dcache__f_reset_reqs__empty_reg )||(! RTL__near_mem__dcache__f_reset_reqs__ENQ && RTL__near_mem__dcache__f_reset_reqs__full_reg ); 
    wire RTL__near_mem__dcache__f_reset_reqs__d1di = RTL__near_mem__dcache__f_reset_reqs__ENQ & RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__f_reset_reqs__CLK )
         begin 
             if ( RTL__near_mem__dcache__f_reset_reqs__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__f_reset_reqs__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__f_reset_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__f_reset_reqs__CLR )
                         begin  
                             RTL__near_mem__dcache__f_reset_reqs__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__f_reset_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__f_reset_reqs__ENQ &&! RTL__near_mem__dcache__f_reset_reqs__DEQ )
                             begin  
                                 RTL__near_mem__dcache__f_reset_reqs__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__f_reset_reqs__full_reg  <=! RTL__near_mem__dcache__f_reset_reqs__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__f_reset_reqs__DEQ &&! RTL__near_mem__dcache__f_reset_reqs__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__f_reset_reqs__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__f_reset_reqs__empty_reg  <=! RTL__near_mem__dcache__f_reset_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__f_reset_reqs__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__f_reset_reqs__data0_reg  <={ RTL__near_mem__dcache__f_reset_reqs__width { RTL__near_mem__dcache__f_reset_reqs__d0di }}& RTL__near_mem__dcache__f_reset_reqs__D_IN |{ RTL__near_mem__dcache__f_reset_reqs__width { RTL__near_mem__dcache__f_reset_reqs__d0d1 }}& RTL__near_mem__dcache__f_reset_reqs__data1_reg |{ RTL__near_mem__dcache__f_reset_reqs__width { RTL__near_mem__dcache__f_reset_reqs__d0h }}& RTL__near_mem__dcache__f_reset_reqs__data0_reg ; 
                 RTL__near_mem__dcache__f_reset_reqs__data1_reg  <= RTL__near_mem__dcache__f_reset_reqs__d1di  ?  RTL__near_mem__dcache__f_reset_reqs__D_IN : RTL__near_mem__dcache__f_reset_reqs__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__f_reset_reqs__CLK )
         begin : RTL__near_mem__dcache__f_reset_reqs__error_checks 
           reg RTL__near_mem__dcache__f_reset_reqs__deqerror , RTL__near_mem__dcache__f_reset_reqs__enqerror ; 
             RTL__near_mem__dcache__f_reset_reqs__deqerror  =0; 
             RTL__near_mem__dcache__f_reset_reqs__enqerror  =0;
             if ( RTL__near_mem__dcache__f_reset_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__f_reset_reqs__empty_reg && RTL__near_mem__dcache__f_reset_reqs__DEQ )
                         begin  
                             RTL__near_mem__dcache__f_reset_reqs__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__f_reset_reqs__full_reg && RTL__near_mem__dcache__f_reset_reqs__ENQ &&(! RTL__near_mem__dcache__f_reset_reqs__DEQ || RTL__near_mem__dcache__f_reset_reqs__guarded ))
                         begin  
                             RTL__near_mem__dcache__f_reset_reqs__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__empty_reg ;
    parameter RTL__near_mem__dcache__f_reset_rsps__width =1; parameter RTL__near_mem__dcache__f_reset_rsps__guarded =1; 
    reg RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
    reg RTL__near_mem__dcache__f_reset_rsps__empty_reg ; reg[ RTL__near_mem__dcache__f_reset_rsps__width -1:0] RTL__near_mem__dcache__f_reset_rsps__data0_reg ; reg[ RTL__near_mem__dcache__f_reset_rsps__width -1:0] RTL__near_mem__dcache__f_reset_rsps__data1_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__FULL_N = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__EMPTY_N = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__D_OUT = RTL__near_mem__dcache__f_reset_rsps__data0_reg ; 
    wire RTL__near_mem__dcache__f_reset_rsps__d0di =( RTL__near_mem__dcache__f_reset_rsps__ENQ &&! RTL__near_mem__dcache__f_reset_rsps__empty_reg )||( RTL__near_mem__dcache__f_reset_rsps__ENQ && RTL__near_mem__dcache__f_reset_rsps__DEQ && RTL__near_mem__dcache__f_reset_rsps__full_reg ); 
    wire RTL__near_mem__dcache__f_reset_rsps__d0d1 = RTL__near_mem__dcache__f_reset_rsps__DEQ &&! RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
    wire RTL__near_mem__dcache__f_reset_rsps__d0h =((! RTL__near_mem__dcache__f_reset_rsps__DEQ )&&(! RTL__near_mem__dcache__f_reset_rsps__ENQ ))||(! RTL__near_mem__dcache__f_reset_rsps__DEQ && RTL__near_mem__dcache__f_reset_rsps__empty_reg )||(! RTL__near_mem__dcache__f_reset_rsps__ENQ && RTL__near_mem__dcache__f_reset_rsps__full_reg ); 
    wire RTL__near_mem__dcache__f_reset_rsps__d1di = RTL__near_mem__dcache__f_reset_rsps__ENQ & RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__f_reset_rsps__CLK )
         begin 
             if ( RTL__near_mem__dcache__f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__f_reset_rsps__CLR )
                         begin  
                             RTL__near_mem__dcache__f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__f_reset_rsps__ENQ &&! RTL__near_mem__dcache__f_reset_rsps__DEQ )
                             begin  
                                 RTL__near_mem__dcache__f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__f_reset_rsps__full_reg  <=! RTL__near_mem__dcache__f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__f_reset_rsps__DEQ &&! RTL__near_mem__dcache__f_reset_rsps__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__f_reset_rsps__empty_reg  <=! RTL__near_mem__dcache__f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__f_reset_rsps__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__f_reset_rsps__data0_reg  <={ RTL__near_mem__dcache__f_reset_rsps__width { RTL__near_mem__dcache__f_reset_rsps__d0di }}& RTL__near_mem__dcache__f_reset_rsps__D_IN |{ RTL__near_mem__dcache__f_reset_rsps__width { RTL__near_mem__dcache__f_reset_rsps__d0d1 }}& RTL__near_mem__dcache__f_reset_rsps__data1_reg |{ RTL__near_mem__dcache__f_reset_rsps__width { RTL__near_mem__dcache__f_reset_rsps__d0h }}& RTL__near_mem__dcache__f_reset_rsps__data0_reg ; 
                 RTL__near_mem__dcache__f_reset_rsps__data1_reg  <= RTL__near_mem__dcache__f_reset_rsps__d1di  ?  RTL__near_mem__dcache__f_reset_rsps__D_IN : RTL__near_mem__dcache__f_reset_rsps__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__f_reset_rsps__CLK )
         begin : RTL__near_mem__dcache__f_reset_rsps__error_checks 
           reg RTL__near_mem__dcache__f_reset_rsps__deqerror , RTL__near_mem__dcache__f_reset_rsps__enqerror ; 
             RTL__near_mem__dcache__f_reset_rsps__deqerror  =0; 
             RTL__near_mem__dcache__f_reset_rsps__enqerror  =0;
             if ( RTL__near_mem__dcache__f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__f_reset_rsps__empty_reg && RTL__near_mem__dcache__f_reset_rsps__DEQ )
                         begin  
                             RTL__near_mem__dcache__f_reset_rsps__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__f_reset_rsps__full_reg && RTL__near_mem__dcache__f_reset_rsps__ENQ &&(! RTL__near_mem__dcache__f_reset_rsps__DEQ || RTL__near_mem__dcache__f_reset_rsps__guarded ))
                         begin  
                             RTL__near_mem__dcache__f_reset_rsps__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__empty_reg ;
    parameter RTL__near_mem__dcache__master_xactor_f_rd_addr__width =1; parameter RTL__near_mem__dcache__master_xactor_f_rd_addr__guarded =1; 
    reg RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
    reg RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_rd_addr__width -1:0] RTL__near_mem__dcache__master_xactor_f_rd_addr__data0_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_rd_addr__width -1:0] RTL__near_mem__dcache__master_xactor_f_rd_addr__data1_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__FULL_N = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__EMPTY_N = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__D_OUT = RTL__near_mem__dcache__master_xactor_f_rd_addr__data0_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__d0di =( RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ &&! RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg )||( RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ && RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ && RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__d0d1 = RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ &&! RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__d0h =((! RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ )&&(! RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ ))||(! RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ && RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg )||(! RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ && RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_rd_addr__d1di = RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ & RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_rd_addr__CLK )
         begin 
             if ( RTL__near_mem__dcache__master_xactor_f_rd_addr__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__master_xactor_f_rd_addr__CLR )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ &&! RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ )
                             begin  
                                 RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg  <=! RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ &&! RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg  <=! RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_rd_addr__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__master_xactor_f_rd_addr__data0_reg  <={ RTL__near_mem__dcache__master_xactor_f_rd_addr__width { RTL__near_mem__dcache__master_xactor_f_rd_addr__d0di }}& RTL__near_mem__dcache__master_xactor_f_rd_addr__D_IN |{ RTL__near_mem__dcache__master_xactor_f_rd_addr__width { RTL__near_mem__dcache__master_xactor_f_rd_addr__d0d1 }}& RTL__near_mem__dcache__master_xactor_f_rd_addr__data1_reg |{ RTL__near_mem__dcache__master_xactor_f_rd_addr__width { RTL__near_mem__dcache__master_xactor_f_rd_addr__d0h }}& RTL__near_mem__dcache__master_xactor_f_rd_addr__data0_reg ; 
                 RTL__near_mem__dcache__master_xactor_f_rd_addr__data1_reg  <= RTL__near_mem__dcache__master_xactor_f_rd_addr__d1di  ?  RTL__near_mem__dcache__master_xactor_f_rd_addr__D_IN : RTL__near_mem__dcache__master_xactor_f_rd_addr__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_rd_addr__CLK )
         begin : RTL__near_mem__dcache__master_xactor_f_rd_addr__error_checks 
           reg RTL__near_mem__dcache__master_xactor_f_rd_addr__deqerror , RTL__near_mem__dcache__master_xactor_f_rd_addr__enqerror ; 
             RTL__near_mem__dcache__master_xactor_f_rd_addr__deqerror  =0; 
             RTL__near_mem__dcache__master_xactor_f_rd_addr__enqerror  =0;
             if ( RTL__near_mem__dcache__master_xactor_f_rd_addr__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg && RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_rd_addr__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg && RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ &&(! RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ || RTL__near_mem__dcache__master_xactor_f_rd_addr__guarded ))
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_rd_addr__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__empty_reg ;
    parameter RTL__near_mem__dcache__master_xactor_f_rd_data__width =1; parameter RTL__near_mem__dcache__master_xactor_f_rd_data__guarded =1; 
    reg RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
    reg RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_rd_data__width -1:0] RTL__near_mem__dcache__master_xactor_f_rd_data__data0_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_rd_data__width -1:0] RTL__near_mem__dcache__master_xactor_f_rd_data__data1_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__FULL_N = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__EMPTY_N = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__D_OUT = RTL__near_mem__dcache__master_xactor_f_rd_data__data0_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__d0di =( RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ &&! RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg )||( RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ && RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ && RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__d0d1 = RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ &&! RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__d0h =((! RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ )&&(! RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ ))||(! RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ && RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg )||(! RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ && RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_rd_data__d1di = RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ & RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_rd_data__CLK )
         begin 
             if ( RTL__near_mem__dcache__master_xactor_f_rd_data__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__master_xactor_f_rd_data__CLR )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ &&! RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ )
                             begin  
                                 RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg  <=! RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ &&! RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg  <=! RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_rd_data__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__master_xactor_f_rd_data__data0_reg  <={ RTL__near_mem__dcache__master_xactor_f_rd_data__width { RTL__near_mem__dcache__master_xactor_f_rd_data__d0di }}& RTL__near_mem__dcache__master_xactor_f_rd_data__D_IN |{ RTL__near_mem__dcache__master_xactor_f_rd_data__width { RTL__near_mem__dcache__master_xactor_f_rd_data__d0d1 }}& RTL__near_mem__dcache__master_xactor_f_rd_data__data1_reg |{ RTL__near_mem__dcache__master_xactor_f_rd_data__width { RTL__near_mem__dcache__master_xactor_f_rd_data__d0h }}& RTL__near_mem__dcache__master_xactor_f_rd_data__data0_reg ; 
                 RTL__near_mem__dcache__master_xactor_f_rd_data__data1_reg  <= RTL__near_mem__dcache__master_xactor_f_rd_data__d1di  ?  RTL__near_mem__dcache__master_xactor_f_rd_data__D_IN : RTL__near_mem__dcache__master_xactor_f_rd_data__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_rd_data__CLK )
         begin : RTL__near_mem__dcache__master_xactor_f_rd_data__error_checks 
           reg RTL__near_mem__dcache__master_xactor_f_rd_data__deqerror , RTL__near_mem__dcache__master_xactor_f_rd_data__enqerror ; 
             RTL__near_mem__dcache__master_xactor_f_rd_data__deqerror  =0; 
             RTL__near_mem__dcache__master_xactor_f_rd_data__enqerror  =0;
             if ( RTL__near_mem__dcache__master_xactor_f_rd_data__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg && RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_rd_data__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg && RTL__near_mem__dcache__master_xactor_f_rd_data__ENQ &&(! RTL__near_mem__dcache__master_xactor_f_rd_data__DEQ || RTL__near_mem__dcache__master_xactor_f_rd_data__guarded ))
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_rd_data__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__empty_reg ;
    parameter RTL__near_mem__dcache__master_xactor_f_wr_addr__width =1; parameter RTL__near_mem__dcache__master_xactor_f_wr_addr__guarded =1; 
    reg RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
    reg RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_wr_addr__width -1:0] RTL__near_mem__dcache__master_xactor_f_wr_addr__data0_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_wr_addr__width -1:0] RTL__near_mem__dcache__master_xactor_f_wr_addr__data1_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__FULL_N = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__EMPTY_N = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__D_OUT = RTL__near_mem__dcache__master_xactor_f_wr_addr__data0_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__d0di =( RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ &&! RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg )||( RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ && RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ && RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__d0d1 = RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ &&! RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__d0h =((! RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ )&&(! RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ ))||(! RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ && RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg )||(! RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ && RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_wr_addr__d1di = RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ & RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_addr__CLK )
         begin 
             if ( RTL__near_mem__dcache__master_xactor_f_wr_addr__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__master_xactor_f_wr_addr__CLR )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ &&! RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ )
                             begin  
                                 RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg  <=! RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ &&! RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg  <=! RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_addr__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__master_xactor_f_wr_addr__data0_reg  <={ RTL__near_mem__dcache__master_xactor_f_wr_addr__width { RTL__near_mem__dcache__master_xactor_f_wr_addr__d0di }}& RTL__near_mem__dcache__master_xactor_f_wr_addr__D_IN |{ RTL__near_mem__dcache__master_xactor_f_wr_addr__width { RTL__near_mem__dcache__master_xactor_f_wr_addr__d0d1 }}& RTL__near_mem__dcache__master_xactor_f_wr_addr__data1_reg |{ RTL__near_mem__dcache__master_xactor_f_wr_addr__width { RTL__near_mem__dcache__master_xactor_f_wr_addr__d0h }}& RTL__near_mem__dcache__master_xactor_f_wr_addr__data0_reg ; 
                 RTL__near_mem__dcache__master_xactor_f_wr_addr__data1_reg  <= RTL__near_mem__dcache__master_xactor_f_wr_addr__d1di  ?  RTL__near_mem__dcache__master_xactor_f_wr_addr__D_IN : RTL__near_mem__dcache__master_xactor_f_wr_addr__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_addr__CLK )
         begin : RTL__near_mem__dcache__master_xactor_f_wr_addr__error_checks 
           reg RTL__near_mem__dcache__master_xactor_f_wr_addr__deqerror , RTL__near_mem__dcache__master_xactor_f_wr_addr__enqerror ; 
             RTL__near_mem__dcache__master_xactor_f_wr_addr__deqerror  =0; 
             RTL__near_mem__dcache__master_xactor_f_wr_addr__enqerror  =0;
             if ( RTL__near_mem__dcache__master_xactor_f_wr_addr__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg && RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_addr__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg && RTL__near_mem__dcache__master_xactor_f_wr_addr__ENQ &&(! RTL__near_mem__dcache__master_xactor_f_wr_addr__DEQ || RTL__near_mem__dcache__master_xactor_f_wr_addr__guarded ))
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_addr__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__empty_reg ;
    parameter RTL__near_mem__dcache__master_xactor_f_wr_data__width =1; parameter RTL__near_mem__dcache__master_xactor_f_wr_data__guarded =1; 
    reg RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
    reg RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_wr_data__width -1:0] RTL__near_mem__dcache__master_xactor_f_wr_data__data0_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_wr_data__width -1:0] RTL__near_mem__dcache__master_xactor_f_wr_data__data1_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__FULL_N = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__EMPTY_N = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__D_OUT = RTL__near_mem__dcache__master_xactor_f_wr_data__data0_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__d0di =( RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ &&! RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg )||( RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ && RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ && RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__d0d1 = RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ &&! RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__d0h =((! RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ )&&(! RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ ))||(! RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ && RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg )||(! RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ && RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_wr_data__d1di = RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ & RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_data__CLK )
         begin 
             if ( RTL__near_mem__dcache__master_xactor_f_wr_data__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__master_xactor_f_wr_data__CLR )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ &&! RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ )
                             begin  
                                 RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg  <=! RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ &&! RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg  <=! RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_data__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__master_xactor_f_wr_data__data0_reg  <={ RTL__near_mem__dcache__master_xactor_f_wr_data__width { RTL__near_mem__dcache__master_xactor_f_wr_data__d0di }}& RTL__near_mem__dcache__master_xactor_f_wr_data__D_IN |{ RTL__near_mem__dcache__master_xactor_f_wr_data__width { RTL__near_mem__dcache__master_xactor_f_wr_data__d0d1 }}& RTL__near_mem__dcache__master_xactor_f_wr_data__data1_reg |{ RTL__near_mem__dcache__master_xactor_f_wr_data__width { RTL__near_mem__dcache__master_xactor_f_wr_data__d0h }}& RTL__near_mem__dcache__master_xactor_f_wr_data__data0_reg ; 
                 RTL__near_mem__dcache__master_xactor_f_wr_data__data1_reg  <= RTL__near_mem__dcache__master_xactor_f_wr_data__d1di  ?  RTL__near_mem__dcache__master_xactor_f_wr_data__D_IN : RTL__near_mem__dcache__master_xactor_f_wr_data__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_data__CLK )
         begin : RTL__near_mem__dcache__master_xactor_f_wr_data__error_checks 
           reg RTL__near_mem__dcache__master_xactor_f_wr_data__deqerror , RTL__near_mem__dcache__master_xactor_f_wr_data__enqerror ; 
             RTL__near_mem__dcache__master_xactor_f_wr_data__deqerror  =0; 
             RTL__near_mem__dcache__master_xactor_f_wr_data__enqerror  =0;
             if ( RTL__near_mem__dcache__master_xactor_f_wr_data__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg && RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_data__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg && RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ &&(! RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ || RTL__near_mem__dcache__master_xactor_f_wr_data__guarded ))
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_data__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__empty_reg ;
    parameter RTL__near_mem__dcache__master_xactor_f_wr_resp__width =1; parameter RTL__near_mem__dcache__master_xactor_f_wr_resp__guarded =1; 
    reg RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
    reg RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_wr_resp__width -1:0] RTL__near_mem__dcache__master_xactor_f_wr_resp__data0_reg ; reg[ RTL__near_mem__dcache__master_xactor_f_wr_resp__width -1:0] RTL__near_mem__dcache__master_xactor_f_wr_resp__data1_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__FULL_N = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__EMPTY_N = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__D_OUT = RTL__near_mem__dcache__master_xactor_f_wr_resp__data0_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__d0di =( RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ &&! RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg )||( RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ && RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ && RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__d0d1 = RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ &&! RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__d0h =((! RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ )&&(! RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ ))||(! RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ && RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg )||(! RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ && RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ); 
    wire RTL__near_mem__dcache__master_xactor_f_wr_resp__d1di = RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ & RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_resp__CLK )
         begin 
             if ( RTL__near_mem__dcache__master_xactor_f_wr_resp__RST ==1'b0)
                 begin  
                     RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg  <=1'b0; 
                     RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__master_xactor_f_wr_resp__CLR )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg  <=1'b0; 
                             RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ &&! RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ )
                             begin  
                                 RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg  <=1'b1; 
                                 RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg  <=! RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ &&! RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ )
                                 begin  
                                     RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg  <=1'b1; 
                                     RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg  <=! RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_resp__CLK )
         begin 
             begin  
                 RTL__near_mem__dcache__master_xactor_f_wr_resp__data0_reg  <={ RTL__near_mem__dcache__master_xactor_f_wr_resp__width { RTL__near_mem__dcache__master_xactor_f_wr_resp__d0di }}& RTL__near_mem__dcache__master_xactor_f_wr_resp__D_IN |{ RTL__near_mem__dcache__master_xactor_f_wr_resp__width { RTL__near_mem__dcache__master_xactor_f_wr_resp__d0d1 }}& RTL__near_mem__dcache__master_xactor_f_wr_resp__data1_reg |{ RTL__near_mem__dcache__master_xactor_f_wr_resp__width { RTL__near_mem__dcache__master_xactor_f_wr_resp__d0h }}& RTL__near_mem__dcache__master_xactor_f_wr_resp__data0_reg ; 
                 RTL__near_mem__dcache__master_xactor_f_wr_resp__data1_reg  <= RTL__near_mem__dcache__master_xactor_f_wr_resp__d1di  ?  RTL__near_mem__dcache__master_xactor_f_wr_resp__D_IN : RTL__near_mem__dcache__master_xactor_f_wr_resp__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__dcache__master_xactor_f_wr_resp__CLK )
         begin : RTL__near_mem__dcache__master_xactor_f_wr_resp__error_checks 
           reg RTL__near_mem__dcache__master_xactor_f_wr_resp__deqerror , RTL__near_mem__dcache__master_xactor_f_wr_resp__enqerror ; 
             RTL__near_mem__dcache__master_xactor_f_wr_resp__deqerror  =0; 
             RTL__near_mem__dcache__master_xactor_f_wr_resp__enqerror  =0;
             if ( RTL__near_mem__dcache__master_xactor_f_wr_resp__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg && RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ )
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_resp__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg && RTL__near_mem__dcache__master_xactor_f_wr_resp__ENQ &&(! RTL__near_mem__dcache__master_xactor_f_wr_resp__DEQ || RTL__near_mem__dcache__master_xactor_f_wr_resp__guarded ))
                         begin  
                             RTL__near_mem__dcache__master_xactor_f_wr_resp__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__empty_reg ;
      
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset__CLKA;
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset__ENA;
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset__WEA;
    wire[RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDR_WIDTH-1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDRA;
    wire[RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DIA;
    wire[RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA;
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset__CLKB;
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset__ENB;
    wire RTL__near_mem__dcache__ram_state_and_ctag_cset__WEB;
    wire[RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDR_WIDTH-1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDRB;
    wire[RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DIB;
    wire[RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB;
    wire RTL__near_mem__dcache__ram_word64_set__CLKA;
    wire RTL__near_mem__dcache__ram_word64_set__ENA;
    wire RTL__near_mem__dcache__ram_word64_set__WEA;
    wire[RTL__near_mem__dcache__ram_word64_set__ADDR_WIDTH-1:0] RTL__near_mem__dcache__ram_word64_set__ADDRA;
    wire[RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_word64_set__DIA;
    wire[RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_word64_set__DOA;
    wire RTL__near_mem__dcache__ram_word64_set__CLKB;
    wire RTL__near_mem__dcache__ram_word64_set__ENB;
    wire RTL__near_mem__dcache__ram_word64_set__WEB;
    wire[RTL__near_mem__dcache__ram_word64_set__ADDR_WIDTH-1:0] RTL__near_mem__dcache__ram_word64_set__ADDRB;
    wire[RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_word64_set__DIB;
    wire[RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__dcache__ram_word64_set__DOB;
    wire RTL__near_mem__icache__ram_state_and_ctag_cset__CLKA;
    wire RTL__near_mem__icache__ram_state_and_ctag_cset__ENA;
    wire RTL__near_mem__icache__ram_state_and_ctag_cset__WEA;
    wire[RTL__near_mem__icache__ram_state_and_ctag_cset__ADDR_WIDTH-1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__ADDRA;
    wire[RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DIA;
    wire[RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DOA;
    wire RTL__near_mem__icache__ram_state_and_ctag_cset__CLKB;
    wire RTL__near_mem__icache__ram_state_and_ctag_cset__ENB;
    wire RTL__near_mem__icache__ram_state_and_ctag_cset__WEB;
    wire[RTL__near_mem__icache__ram_state_and_ctag_cset__ADDR_WIDTH-1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__ADDRB;
    wire[RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DIB;
    wire[RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DOB;
    wire RTL__near_mem__icache__ram_word64_set__CLKA;
    wire RTL__near_mem__icache__ram_word64_set__ENA;
    wire RTL__near_mem__icache__ram_word64_set__WEA;
    wire[RTL__near_mem__icache__ram_word64_set__ADDR_WIDTH-1:0] RTL__near_mem__icache__ram_word64_set__ADDRA;
    wire[RTL__near_mem__icache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_word64_set__DIA;
    wire[RTL__near_mem__icache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_word64_set__DOA;
    wire RTL__near_mem__icache__ram_word64_set__CLKB;
    wire RTL__near_mem__icache__ram_word64_set__ENB;
    wire RTL__near_mem__icache__ram_word64_set__WEB;
    wire[RTL__near_mem__icache__ram_word64_set__ADDR_WIDTH-1:0] RTL__near_mem__icache__ram_word64_set__ADDRB;
    wire[RTL__near_mem__icache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_word64_set__DIB;
    wire[RTL__near_mem__icache__ram_word64_set__DATA_WIDTH-1:0] RTL__near_mem__icache__ram_word64_set__DOB;

    reg[ RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R ; reg[ RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R ; reg[ RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R2 ; reg[ RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R2 ; parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__PIPELINED =0; parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDR_WIDTH =1; parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH =1; parameter RTL__near_mem__dcache__ram_state_and_ctag_cset__MEMSIZE =1; (* RTL__near_mem__dcache__ram_state_and_ctag_cset__keep *)
    wire[ RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__arb1 ; (* RTL__near_mem__dcache__ram_state_and_ctag_cset__keep *)
    wire[ RTL__near_mem__dcache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_state_and_ctag_cset__arb2 ; 
  always @( posedge  RTL__near_mem__dcache__ram_state_and_ctag_cset__CLKA )
         begin 
             if ( RTL__near_mem__dcache__ram_state_and_ctag_cset__ENA )
                 begin 
                     if ( RTL__near_mem__dcache__ram_state_and_ctag_cset__WEA )
                         begin  
                             RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R  <= RTL__near_mem__dcache__ram_state_and_ctag_cset__DIA ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R  <= RTL__near_mem__dcache__ram_state_and_ctag_cset__arb1 ;
                         end 
                 end  
             RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R2  <= RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R ;
         end
  always @( posedge  RTL__near_mem__dcache__ram_state_and_ctag_cset__CLKB )
         begin 
             if ( RTL__near_mem__dcache__ram_state_and_ctag_cset__ENB )
                 begin 
                     if ( RTL__near_mem__dcache__ram_state_and_ctag_cset__WEB )
                         begin  
                             RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R  <= RTL__near_mem__dcache__ram_state_and_ctag_cset__DIB ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R  <= RTL__near_mem__dcache__ram_state_and_ctag_cset__arb2 ;
                         end 
                 end  
             RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R2  <= RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R ;
         end
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA =( RTL__near_mem__dcache__ram_state_and_ctag_cset__PIPELINED ) ?  RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R2 : RTL__near_mem__dcache__ram_state_and_ctag_cset__DOA_R ; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB =( RTL__near_mem__dcache__ram_state_and_ctag_cset__PIPELINED ) ?  RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R2 : RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB_R ;
    reg[ RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_word64_set__DOA_R ; reg[ RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_word64_set__DOB_R ; reg[ RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_word64_set__DOA_R2 ; reg[ RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_word64_set__DOB_R2 ; parameter RTL__near_mem__dcache__ram_word64_set__PIPELINED =0; parameter RTL__near_mem__dcache__ram_word64_set__ADDR_WIDTH =1; parameter RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH =1; parameter RTL__near_mem__dcache__ram_word64_set__MEMSIZE =1; (* RTL__near_mem__dcache__ram_word64_set__keep *)
    wire[ RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_word64_set__arb1 ; (* RTL__near_mem__dcache__ram_word64_set__keep *)
    wire[ RTL__near_mem__dcache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__dcache__ram_word64_set__arb2 ; 
  always @( posedge  RTL__near_mem__dcache__ram_word64_set__CLKA )
         begin 
             if ( RTL__near_mem__dcache__ram_word64_set__ENA )
                 begin 
                     if ( RTL__near_mem__dcache__ram_word64_set__WEA )
                         begin  
                             RTL__near_mem__dcache__ram_word64_set__DOA_R  <= RTL__near_mem__dcache__ram_word64_set__DIA ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__dcache__ram_word64_set__DOA_R  <= RTL__near_mem__dcache__ram_word64_set__arb1 ;
                         end 
                 end  
             RTL__near_mem__dcache__ram_word64_set__DOA_R2  <= RTL__near_mem__dcache__ram_word64_set__DOA_R ;
         end
  always @( posedge  RTL__near_mem__dcache__ram_word64_set__CLKB )
         begin 
             if ( RTL__near_mem__dcache__ram_word64_set__ENB )
                 begin 
                     if ( RTL__near_mem__dcache__ram_word64_set__WEB )
                         begin  
                             RTL__near_mem__dcache__ram_word64_set__DOB_R  <= RTL__near_mem__dcache__ram_word64_set__DIB ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__dcache__ram_word64_set__DOB_R  <= RTL__near_mem__dcache__ram_word64_set__arb2 ;
                         end 
                 end  
             RTL__near_mem__dcache__ram_word64_set__DOB_R2  <= RTL__near_mem__dcache__ram_word64_set__DOB_R ;
         end
  assign  RTL__near_mem__dcache__ram_word64_set__DOA =( RTL__near_mem__dcache__ram_word64_set__PIPELINED ) ?  RTL__near_mem__dcache__ram_word64_set__DOA_R2 : RTL__near_mem__dcache__ram_word64_set__DOA_R ; 
  assign  RTL__near_mem__dcache__ram_word64_set__DOB =( RTL__near_mem__dcache__ram_word64_set__PIPELINED ) ?  RTL__near_mem__dcache__ram_word64_set__DOB_R2 : RTL__near_mem__dcache__ram_word64_set__DOB_R ;
      
    wire RTL__near_mem__dcache__soc_map__CLK;
    wire RTL__near_mem__dcache__soc_map__RST_N;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_base;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_size;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_lim;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_plic_addr_base;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_plic_addr_size;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_plic_addr_lim;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_uart0_addr_base;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_uart0_addr_size;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_uart0_addr_lim;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_boot_rom_addr_base;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_boot_rom_addr_size;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_boot_rom_addr_lim;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_base;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_size;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_lim;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_tcm_addr_base;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_tcm_addr_size;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_tcm_addr_lim;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_is_mem_addr_addr;
    wire RTL__near_mem__dcache__soc_map__m_is_mem_addr;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr;
    wire RTL__near_mem__dcache__soc_map__m_is_IO_addr;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr_addr;
    wire RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_pc_reset_value;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_mtvec_reset_value;
    wire[63:0] RTL__near_mem__dcache__soc_map__m_nmivec_reset_value;
    wire RTL__near_mem__icache__soc_map__CLK;
    wire RTL__near_mem__icache__soc_map__RST_N;
    wire[63:0] RTL__near_mem__icache__soc_map__m_near_mem_io_addr_base;
    wire[63:0] RTL__near_mem__icache__soc_map__m_near_mem_io_addr_size;
    wire[63:0] RTL__near_mem__icache__soc_map__m_near_mem_io_addr_lim;
    wire[63:0] RTL__near_mem__icache__soc_map__m_plic_addr_base;
    wire[63:0] RTL__near_mem__icache__soc_map__m_plic_addr_size;
    wire[63:0] RTL__near_mem__icache__soc_map__m_plic_addr_lim;
    wire[63:0] RTL__near_mem__icache__soc_map__m_uart0_addr_base;
    wire[63:0] RTL__near_mem__icache__soc_map__m_uart0_addr_size;
    wire[63:0] RTL__near_mem__icache__soc_map__m_uart0_addr_lim;
    wire[63:0] RTL__near_mem__icache__soc_map__m_boot_rom_addr_base;
    wire[63:0] RTL__near_mem__icache__soc_map__m_boot_rom_addr_size;
    wire[63:0] RTL__near_mem__icache__soc_map__m_boot_rom_addr_lim;
    wire[63:0] RTL__near_mem__icache__soc_map__m_mem0_controller_addr_base;
    wire[63:0] RTL__near_mem__icache__soc_map__m_mem0_controller_addr_size;
    wire[63:0] RTL__near_mem__icache__soc_map__m_mem0_controller_addr_lim;
    wire[63:0] RTL__near_mem__icache__soc_map__m_tcm_addr_base;
    wire[63:0] RTL__near_mem__icache__soc_map__m_tcm_addr_size;
    wire[63:0] RTL__near_mem__icache__soc_map__m_tcm_addr_lim;
    wire[63:0] RTL__near_mem__icache__soc_map__m_is_mem_addr_addr;
    wire RTL__near_mem__icache__soc_map__m_is_mem_addr;
    wire[63:0] RTL__near_mem__icache__soc_map__m_is_IO_addr_addr;
    wire RTL__near_mem__icache__soc_map__m_is_IO_addr;
    wire[63:0] RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr_addr;
    wire RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr;
    wire[63:0] RTL__near_mem__icache__soc_map__m_pc_reset_value;
    wire[63:0] RTL__near_mem__icache__soc_map__m_mtvec_reset_value;
    wire[63:0] RTL__near_mem__icache__soc_map__m_nmivec_reset_value;
    wire RTL__near_mem__soc_map__CLK;
    wire RTL__near_mem__soc_map__RST_N;
    wire[63:0] RTL__near_mem__soc_map__m_near_mem_io_addr_base;
    wire[63:0] RTL__near_mem__soc_map__m_near_mem_io_addr_size;
    wire[63:0] RTL__near_mem__soc_map__m_near_mem_io_addr_lim;
    wire[63:0] RTL__near_mem__soc_map__m_plic_addr_base;
    wire[63:0] RTL__near_mem__soc_map__m_plic_addr_size;
    wire[63:0] RTL__near_mem__soc_map__m_plic_addr_lim;
    wire[63:0] RTL__near_mem__soc_map__m_uart0_addr_base;
    wire[63:0] RTL__near_mem__soc_map__m_uart0_addr_size;
    wire[63:0] RTL__near_mem__soc_map__m_uart0_addr_lim;
    wire[63:0] RTL__near_mem__soc_map__m_boot_rom_addr_base;
    wire[63:0] RTL__near_mem__soc_map__m_boot_rom_addr_size;
    wire[63:0] RTL__near_mem__soc_map__m_boot_rom_addr_lim;
    wire[63:0] RTL__near_mem__soc_map__m_mem0_controller_addr_base;
    wire[63:0] RTL__near_mem__soc_map__m_mem0_controller_addr_size;
    wire[63:0] RTL__near_mem__soc_map__m_mem0_controller_addr_lim;
    wire[63:0] RTL__near_mem__soc_map__m_tcm_addr_base;
    wire[63:0] RTL__near_mem__soc_map__m_tcm_addr_size;
    wire[63:0] RTL__near_mem__soc_map__m_tcm_addr_lim;
    wire[63:0] RTL__near_mem__soc_map__m_is_mem_addr_addr;
    wire RTL__near_mem__soc_map__m_is_mem_addr;
    wire[63:0] RTL__near_mem__soc_map__m_is_IO_addr_addr;
    wire RTL__near_mem__soc_map__m_is_IO_addr;
    wire[63:0] RTL__near_mem__soc_map__m_is_near_mem_IO_addr_addr;
    wire RTL__near_mem__soc_map__m_is_near_mem_IO_addr;
    wire[63:0] RTL__near_mem__soc_map__m_pc_reset_value;
    wire[63:0] RTL__near_mem__soc_map__m_mtvec_reset_value;
    wire[63:0] RTL__near_mem__soc_map__m_nmivec_reset_value;

    wire[63:0] RTL__near_mem__dcache__soc_map__m_boot_rom_addr_base , RTL__near_mem__dcache__soc_map__m_boot_rom_addr_lim , RTL__near_mem__dcache__soc_map__m_boot_rom_addr_size , RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_base , RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_lim , RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_size , RTL__near_mem__dcache__soc_map__m_mtvec_reset_value , RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_base , RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_lim , RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_size , RTL__near_mem__dcache__soc_map__m_nmivec_reset_value , RTL__near_mem__dcache__soc_map__m_pc_reset_value , RTL__near_mem__dcache__soc_map__m_plic_addr_base , RTL__near_mem__dcache__soc_map__m_plic_addr_lim , RTL__near_mem__dcache__soc_map__m_plic_addr_size , RTL__near_mem__dcache__soc_map__m_tcm_addr_base , RTL__near_mem__dcache__soc_map__m_tcm_addr_lim , RTL__near_mem__dcache__soc_map__m_tcm_addr_size , RTL__near_mem__dcache__soc_map__m_uart0_addr_base , RTL__near_mem__dcache__soc_map__m_uart0_addr_lim , RTL__near_mem__dcache__soc_map__m_uart0_addr_size ; 
    wire RTL__near_mem__dcache__soc_map__m_is_IO_addr , RTL__near_mem__dcache__soc_map__m_is_mem_addr , RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr ; 
  assign  RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL__near_mem__dcache__soc_map__m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL__near_mem__dcache__soc_map__m_plic_addr_base =64'h000000000C000000; 
  assign  RTL__near_mem__dcache__soc_map__m_plic_addr_size =64'h0000000000400000; 
  assign  RTL__near_mem__dcache__soc_map__m_plic_addr_lim =64'd205520896; 
  assign  RTL__near_mem__dcache__soc_map__m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL__near_mem__dcache__soc_map__m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL__near_mem__dcache__soc_map__m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL__near_mem__dcache__soc_map__m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL__near_mem__dcache__soc_map__m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL__near_mem__dcache__soc_map__m_boot_rom_addr_lim =64'd8192; 
  assign  RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL__near_mem__dcache__soc_map__m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL__near_mem__dcache__soc_map__m_tcm_addr_base =64'h0; 
  assign  RTL__near_mem__dcache__soc_map__m_tcm_addr_size =64'd0; 
  assign  RTL__near_mem__dcache__soc_map__m_tcm_addr_lim =64'd0; 
  assign  RTL__near_mem__dcache__soc_map__m_is_mem_addr = RTL__near_mem__dcache__soc_map__m_is_mem_addr_addr >=64'h0000000000001000&& RTL__near_mem__dcache__soc_map__m_is_mem_addr_addr <64'd8192|| RTL__near_mem__dcache__soc_map__m_is_mem_addr_addr >=64'h0000000080000000&& RTL__near_mem__dcache__soc_map__m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL__near_mem__dcache__soc_map__m_is_IO_addr = RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr >=64'h0000000002000000&& RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr <64'd33603584|| RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr >=64'h000000000C000000&& RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr <64'd205520896|| RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr >=64'h00000000C0000000&& RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr = RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL__near_mem__dcache__soc_map__m_pc_reset_value =64'h0000000000001000; 
  assign  RTL__near_mem__dcache__soc_map__m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL__near_mem__dcache__soc_map__m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
     
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req = RTL__near_mem__dcache__f_fabric_write_reqs$EMPTY_N && RTL__near_mem__dcache__master_xactor_f_wr_addr$FULL_N && RTL__near_mem__dcache__master_xactor_f_wr_data$FULL_N ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req = RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_reset =( RTL__near_mem__dcache__rg_cset_in_cache !=7'd127|| RTL__near_mem__dcache__f_reset_reqs$EMPTY_N && RTL__near_mem__dcache__f_reset_rsps$FULL_N )&& RTL__near_mem__dcache__rg_state ==4'd1; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset = RTL__near_mem__dcache__CAN_FIRE_RL_rl_reset ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_probe_and_immed_rsp =( RTL__near_mem__dcache__dmem_not_imem &&! RTL__near_mem__dcache__soc_map$m_is_mem_addr ||! RTL__near_mem__dcache__rg_op || RTL__near_mem__dcache__f_fabric_write_reqs$FULL_N )&& RTL__near_mem__dcache__rg_state ==4'd3; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp = RTL__near_mem__dcache__CAN_FIRE_RL_rl_probe_and_immed_rsp &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_start_cache_refill = RTL__near_mem__dcache__master_xactor_f_rd_addr$FULL_N && RTL__near_mem__dcache__rg_state ==4'd8&& RTL__near_mem__dcache__b__h14485 ==4'd0; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill = RTL__near_mem__dcache__CAN_FIRE_RL_rl_start_cache_refill &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__EN_req ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_cache_refill_rsps_loop = RTL__near_mem__dcache__master_xactor_f_rd_data$EMPTY_N && RTL__near_mem__dcache__rg_state ==4'd9; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop = RTL__near_mem__dcache__CAN_FIRE_RL_rl_cache_refill_rsps_loop &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__EN_req ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_rereq = RTL__near_mem__dcache__rg_state ==4'd10; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq = RTL__near_mem__dcache__CAN_FIRE_RL_rl_rereq &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__EN_req ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_ST_AMO_response = RTL__near_mem__dcache__rg_state ==4'd11; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_ST_AMO_response = RTL__near_mem__dcache__CAN_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_read_req = RTL__near_mem__dcache__master_xactor_f_rd_addr$FULL_N && RTL__near_mem__dcache__rg_state ==4'd12&&! RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__b__h14485 ==4'd0; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req = RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_read_req &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_read_rsp = RTL__near_mem__dcache__master_xactor_f_rd_data$EMPTY_N && RTL__near_mem__dcache__rg_state ==4'd13; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp = RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_read_rsp &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_maintain_io_read_rsp = RTL__near_mem__dcache__rg_state ==4'd14; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_maintain_io_read_rsp = RTL__near_mem__dcache__CAN_FIRE_RL_rl_maintain_io_read_rsp ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_write_req = RTL__near_mem__dcache__f_fabric_write_reqs$FULL_N && RTL__near_mem__dcache__rg_state ==4'd12&& RTL__near_mem__dcache__rg_op ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req = RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_discard_write_rsp = RTL__near_mem__dcache__b__h14485 !=4'd0&& RTL__near_mem__dcache__master_xactor_f_wr_resp$EMPTY_N ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp = RTL__near_mem__dcache__CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_drive_exception_rsp = RTL__near_mem__dcache__rg_state ==4'd4; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_drive_exception_rsp = RTL__near_mem__dcache__rg_state ==4'd4; 
  assign  RTL__near_mem__dcache__CAN_FIRE_RL_rl_start_reset = RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset = RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_1 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_2 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 ; 
  assign  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__SEL_3 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL__near_mem__dcache__WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__SEL_1 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op ; 
  assign  RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 = RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 ; 
  assign  RTL__near_mem__dcache__MUX_ram_word64_set$a_put_1__SEL_1 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]!=2'd3; 
  assign  RTL__near_mem__dcache__MUX_rg_error_during_refill$write_1__SEL_1 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_1 = RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_2 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_2 = RTL__near_mem__dcache__f_reset_reqs$EMPTY_N && RTL__near_mem__dcache__rg_state !=4'd1; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_3 = RTL__near_mem__dcache__CAN_FIRE_RL_rl_io_write_req &&! RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_7 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]==2'd3; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_9 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 ; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_10 = RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127; 
  always @(          RTL__near_mem__dcache__rg_f3                          or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247                 or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276                or   RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32               or   RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__word64__h5094             or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264            or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285           or   RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  )
         begin 
             case ( RTL__near_mem__dcache__rg_f3 )
              3 'b0: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 ;
              3 'b001: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 ;
              3 'b010: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 ;
              3 'b011: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  =( RTL__near_mem__dcache__rg_addr [2:0]==3'h0) ?  RTL__near_mem__dcache__word64__h5094 :64'd0;
              3 'b100: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 ;
              3 'b101: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 ;
              3 'b110: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 ;
              3 'd7: 
                  RTL__near_mem__dcache__MUX_dw_output_ld_val$wset_1__VAL_2  =64'd0;endcase
         end
  assign  RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__VAL_1 ={ RTL__near_mem__dcache__rg_f3 , RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_st_amo_val }; 
  assign  RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__VAL_2 ={ RTL__near_mem__dcache__rg_f3 , RTL__near_mem__dcache__rg_pa , RTL__near_mem__dcache__rg_st_amo_val }; 
  assign  RTL__near_mem__dcache__MUX_master_xactor_f_rd_addr$enq_1__VAL_1 ={4'd0, RTL__near_mem__dcache__cline_fabric_addr__h14584 ,29'd7143424}; 
  assign  RTL__near_mem__dcache__MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ={4'd0, RTL__near_mem__dcache__fabric_addr__h17243 ,8'd0, RTL__near_mem__dcache__value__h17372 ,18'd65536}; 
  assign  RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ={3'd4, RTL__near_mem__dcache__rg_pa [31:12]}; 
  assign  RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_2 = RTL__near_mem__dcache__rg_word64_set_in_cache +9'd1; 
  assign  RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_4 ={ RTL__near_mem__dcache__rg_addr [11:5],2'd0}; 
  assign  RTL__near_mem__dcache__MUX_rg_cset_in_cache$write_1__VAL_1 = RTL__near_mem__dcache__rg_cset_in_cache +7'd1; 
  assign  RTL__near_mem__dcache__MUX_rg_exc_code$write_1__VAL_1 = RTL__near_mem__dcache__req_op  ? 4'd6:4'd4; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_1 = RTL__near_mem__dcache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539  ? 4'd4:4'd3; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_4 =( RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0) ? 4'd14:4'd4; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_7 =( RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__dcache__rg_error_during_refill ) ? 4'd4:4'd10; 
  assign  RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_9 =( RTL__near_mem__dcache__dmem_not_imem &&! RTL__near_mem__dcache__soc_map$m_is_mem_addr ) ? 4'd12:( RTL__near_mem__dcache__rg_op  ? 4'd11:4'd8); 
  assign  RTL__near_mem__dcache__dw_valid$whas = RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 || RTL__near_mem__dcache__WILL_FIRE_RL_rl_drive_exception_rsp || RTL__near_mem__dcache__WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL__near_mem__dcache__WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port0__write_1 = RTL__near_mem__dcache__ctr_wr_rsps_pending_crg +4'd1; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port1__write_1 = RTL__near_mem__dcache__b__h14485 -4'd1; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port2__read = RTL__near_mem__dcache__CAN_FIRE_RL_rl_discard_write_rsp  ?  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port1__write_1 : RTL__near_mem__dcache__b__h14485 ; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$EN_port2__write = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port3__read = RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$EN_port2__write  ? 4'd0: RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port2__read ; 
  assign  RTL__near_mem__dcache__cfg_verbosity$D_IN = RTL__near_mem__dcache__set_verbosity_verbosity ; 
  assign  RTL__near_mem__dcache__cfg_verbosity$EN = RTL__near_mem__dcache__EN_set_verbosity ; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$D_IN = RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port3__read ; 
  assign  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$EN =1'b1; 
  assign  RTL__near_mem__dcache__rg_addr$D_IN = RTL__near_mem__dcache__req_addr ; 
  assign  RTL__near_mem__dcache__rg_addr$EN = RTL__near_mem__dcache__EN_req ; (* RTL__near_mem__dcache__keep *)
    wire[6:0] RTL__near_mem__dcache__MUX_rg_cset_in_cache$write_1__VAL_1_any_val ; 
  assign  RTL__near_mem__dcache__rg_cset_in_cache$D_IN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset  ?  RTL__near_mem__dcache__MUX_rg_cset_in_cache$write_1__VAL_1_any_val :7'd0; 
  assign  RTL__near_mem__dcache__rg_cset_in_cache$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset || RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__dcache__rg_error_during_refill$D_IN = RTL__near_mem__dcache__MUX_rg_error_during_refill$write_1__SEL_1 ; 
  assign  RTL__near_mem__dcache__rg_error_during_refill$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill ; 
  always @(      RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_1                  or   RTL__near_mem__dcache__MUX_rg_exc_code$write_1__VAL_1             or   RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_2            or   RTL__near_mem__dcache__MUX_rg_error_during_refill$write_1__SEL_1           or   RTL__near_mem__dcache__access_exc_code__h2256  )
         case (1'b1) 
          RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_1  : 
              RTL__near_mem__dcache__rg_exc_code$D_IN  = RTL__near_mem__dcache__MUX_rg_exc_code$write_1__VAL_1 ; 
          RTL__near_mem__dcache__MUX_rg_exc_code$write_1__SEL_2  : 
              RTL__near_mem__dcache__rg_exc_code$D_IN  =4'd5; 
          RTL__near_mem__dcache__MUX_rg_error_during_refill$write_1__SEL_1  : 
              RTL__near_mem__dcache__rg_exc_code$D_IN  = RTL__near_mem__dcache__access_exc_code__h2256 ;
          default : 
              RTL__near_mem__dcache__rg_exc_code$D_IN  =4'b1010;endcase
  assign  RTL__near_mem__dcache__rg_exc_code$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL__near_mem__dcache__rg_f3$D_IN = RTL__near_mem__dcache__req_f3 ; 
  assign  RTL__near_mem__dcache__rg_f3$EN = RTL__near_mem__dcache__EN_req ; 
  assign  RTL__near_mem__dcache__rg_ld_val$D_IN = RTL__near_mem__dcache__ld_val__h17594 ; 
  assign  RTL__near_mem__dcache__rg_ld_val$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp ; 
  assign  RTL__near_mem__dcache__rg_lower_word32$D_IN =32'h0; 
  assign  RTL__near_mem__dcache__rg_lower_word32$EN =1'b0; 
  assign  RTL__near_mem__dcache__rg_lower_word32_full$D_IN =1'd0; 
  assign  RTL__near_mem__dcache__rg_lower_word32_full$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__dcache__rg_op$D_IN = RTL__near_mem__dcache__req_op ; 
  assign  RTL__near_mem__dcache__rg_op$EN = RTL__near_mem__dcache__EN_req ; 
  assign  RTL__near_mem__dcache__rg_pa$D_IN = RTL__near_mem__dcache__EN_req  ?  RTL__near_mem__dcache__req_addr : RTL__near_mem__dcache__rg_addr ; 
  assign  RTL__near_mem__dcache__rg_pa$EN = RTL__near_mem__dcache__EN_req || RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp ; 
  assign  RTL__near_mem__dcache__rg_pte_pa$D_IN =32'h0; 
  assign  RTL__near_mem__dcache__rg_pte_pa$EN =1'b0; 
  assign  RTL__near_mem__dcache__rg_st_amo_val$D_IN = RTL__near_mem__dcache__req_st_value ; 
  assign  RTL__near_mem__dcache__rg_st_amo_val$EN = RTL__near_mem__dcache__EN_req ; 
  always @(               RTL__near_mem__dcache__EN_req                                    or   RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_1                      or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset                     or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req                    or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp                   or   RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_4                  or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req                 or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq                or   RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_7               or   RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_7              or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill             or   RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_9            or   RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_9           or   RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_10  )
         case (1'b1) 
          RTL__near_mem__dcache__EN_req  : 
              RTL__near_mem__dcache__rg_state$D_IN  = RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_1 ; 
          RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset  : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'd1; 
          RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req  : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'd11; 
          RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp  : 
              RTL__near_mem__dcache__rg_state$D_IN  = RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_4 ; 
          RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req  : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'd13; 
          RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq  : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'd3; 
          RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_7  : 
              RTL__near_mem__dcache__rg_state$D_IN  = RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_7 ; 
          RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'd9; 
          RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_9  : 
              RTL__near_mem__dcache__rg_state$D_IN  = RTL__near_mem__dcache__MUX_rg_state$write_1__VAL_9 ; 
          RTL__near_mem__dcache__MUX_rg_state$write_1__SEL_10  : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'd2;
          default : 
              RTL__near_mem__dcache__rg_state$D_IN  =4'b1010;endcase
  assign  RTL__near_mem__dcache__rg_state$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]==2'd3|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 || RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp || RTL__near_mem__dcache__EN_req || RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset || RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq || RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req || RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL__near_mem__dcache__rg_word64_set_in_cache$D_IN = RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2  ?  RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_2 : RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_4 ; 
  assign  RTL__near_mem__dcache__rg_word64_set_in_cache$EN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]!=2'd3|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs$D_IN = RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__SEL_1  ?  RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__VAL_1 : RTL__near_mem__dcache__MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs$ENQ = RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op || RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs$DEQ = RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__dcache__f_fabric_write_reqs$CLR =1'b0; 
  assign  RTL__near_mem__dcache__f_reset_reqs$D_IN =! RTL__near_mem__dcache__EN_server_reset_request_put ; 
  assign  RTL__near_mem__dcache__f_reset_reqs$ENQ = RTL__near_mem__dcache__EN_server_reset_request_put || RTL__near_mem__dcache__EN_server_flush_request_put ; 
  assign  RTL__near_mem__dcache__f_reset_reqs$DEQ = RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127; 
  assign  RTL__near_mem__dcache__f_reset_reqs$CLR =1'b0; 
  assign  RTL__near_mem__dcache__f_reset_rsps$D_IN = RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__f_reset_rsps$ENQ = RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127; 
  assign  RTL__near_mem__dcache__f_reset_rsps$DEQ = RTL__near_mem__dcache__EN_server_flush_response_get || RTL__near_mem__dcache__EN_server_reset_response_get ; 
  assign  RTL__near_mem__dcache__f_reset_rsps$CLR =1'b0; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr$D_IN = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  ?  RTL__near_mem__dcache__MUX_master_xactor_f_rd_addr$enq_1__VAL_1 : RTL__near_mem__dcache__MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr$ENQ = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr$DEQ = RTL__near_mem__dcache__master_xactor_f_rd_addr$EMPTY_N && RTL__near_mem__dcache__mem_master_arready ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_addr$CLR = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data$D_IN ={ RTL__near_mem__dcache__mem_master_rid , RTL__near_mem__dcache__mem_master_rdata , RTL__near_mem__dcache__mem_master_rresp , RTL__near_mem__dcache__mem_master_rlast }; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data$ENQ = RTL__near_mem__dcache__mem_master_rvalid && RTL__near_mem__dcache__master_xactor_f_rd_data$FULL_N ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data$DEQ = RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp || RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop ; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_data$CLR = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr$D_IN ={4'd0, RTL__near_mem__dcache__mem_req_wr_addr_awaddr__h2473 ,8'd0, RTL__near_mem__dcache__x__h2520 ,18'd65536}; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr$ENQ = RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr$DEQ = RTL__near_mem__dcache__master_xactor_f_wr_addr$EMPTY_N && RTL__near_mem__dcache__mem_master_awready ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_addr$CLR = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data$D_IN ={ RTL__near_mem__dcache__mem_req_wr_data_wdata__h2699 , RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700 ,1'd1}; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data$ENQ = RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data$DEQ = RTL__near_mem__dcache__master_xactor_f_wr_data$EMPTY_N && RTL__near_mem__dcache__mem_master_wready ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_data$CLR = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp$D_IN ={ RTL__near_mem__dcache__mem_master_bid , RTL__near_mem__dcache__mem_master_bresp }; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp$ENQ = RTL__near_mem__dcache__mem_master_bvalid && RTL__near_mem__dcache__master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp$DEQ = RTL__near_mem__dcache__CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL__near_mem__dcache__master_xactor_f_wr_resp$CLR = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__dcache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$ADDRA = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  ?  RTL__near_mem__dcache__rg_addr [11:5]: RTL__near_mem__dcache__rg_cset_in_cache ; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$ADDRB = RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ?  RTL__near_mem__dcache__req_addr [11:5]: RTL__near_mem__dcache__rg_addr [11:5]; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$DIA = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  ?  RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 :23'd2796202; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$DIB = RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ? 23'b01010101010101010101010:23'b01010101010101010101010; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$WEA =1'd1; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$WEB =1'd0; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$ENA = RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset ; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset$ENB = RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq ; 
  assign  RTL__near_mem__dcache__ram_word64_set$ADDRA = RTL__near_mem__dcache__MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL__near_mem__dcache__rg_word64_set_in_cache : RTL__near_mem__dcache__rg_addr [11:3]; 
  always @(         RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                        or   RTL__near_mem__dcache__req_addr                or   RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2               or   RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_2              or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq             or   RTL__near_mem__dcache__rg_addr            or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill           or   RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_4  )
         begin 
             case (1'b1) 
              RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL__near_mem__dcache__ram_word64_set$ADDRB  = RTL__near_mem__dcache__req_addr [11:3]; 
              RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL__near_mem__dcache__ram_word64_set$ADDRB  = RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_2 ; 
              RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq  : 
                  RTL__near_mem__dcache__ram_word64_set$ADDRB  = RTL__near_mem__dcache__rg_addr [11:3]; 
              RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL__near_mem__dcache__ram_word64_set$ADDRB  = RTL__near_mem__dcache__MUX_ram_word64_set$b_put_2__VAL_4 ;
              default : 
                  RTL__near_mem__dcache__ram_word64_set$ADDRB  =9'b010101010;endcase
         end
  assign  RTL__near_mem__dcache__ram_word64_set$DIA = RTL__near_mem__dcache__MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:3]: RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 ; 
  always @(     RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                or   RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2            or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq           or   RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  )
         begin 
             case (1'b1) 
              RTL__near_mem__dcache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL__near_mem__dcache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL__near_mem__dcache__MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL__near_mem__dcache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq  : 
                  RTL__near_mem__dcache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL__near_mem__dcache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;
              default : 
                  RTL__near_mem__dcache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL__near_mem__dcache__ram_word64_set$WEA =1'd1; 
  assign  RTL__near_mem__dcache__ram_word64_set$WEB =1'd0; 
  assign  RTL__near_mem__dcache__ram_word64_set$ENA = RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 ; 
  assign  RTL__near_mem__dcache__ram_word64_set$ENB = RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]!=2'd3|| RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq || RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL__near_mem__dcache__soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL__near_mem__dcache__soc_map$m_is_mem_addr_addr ={32'd0, RTL__near_mem__dcache__rg_addr }; 
  assign  RTL__near_mem__dcache__soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 = RTL__near_mem__dcache__cfg_verbosity >4'd1; 
  assign  RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 = RTL__near_mem__dcache__cfg_verbosity >4'd2; 
  assign  RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 =(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL__near_mem__dcache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 =(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&&! RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL__near_mem__dcache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 = RTL__near_mem__dcache__req_f3 [1:0]!=2'b0&&( RTL__near_mem__dcache__req_f3 [1:0]!=2'b01|| RTL__near_mem__dcache__req_addr [0])&&( RTL__near_mem__dcache__req_f3 [1:0]!=2'b10|| RTL__near_mem__dcache__req_addr [1:0]!=2'b0)&&( RTL__near_mem__dcache__req_f3 [1:0]!=2'b11|| RTL__near_mem__dcache__req_addr [2:0]!=3'b0); 
  assign  RTL__near_mem__dcache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 =! RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL__near_mem__dcache___theResult___snd_fst__h2707 = RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [63:0]<< RTL__near_mem__dcache__shift_bits__h2487 ; 
  assign  RTL__near_mem__dcache__access_exc_code__h2256 = RTL__near_mem__dcache__dmem_not_imem  ? ( RTL__near_mem__dcache__rg_op  ? 4'd7:4'd5):4'd1; 
  assign  RTL__near_mem__dcache__b__h14485 = RTL__near_mem__dcache__CAN_FIRE_RL_rl_fabric_send_write_req  ?  RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$port0__write_1 : RTL__near_mem__dcache__ctr_wr_rsps_pending_crg ; 
  assign  RTL__near_mem__dcache__cline_addr__h14583 ={ RTL__near_mem__dcache__rg_pa [31:5],5'd0}; 
  assign  RTL__near_mem__dcache__cline_fabric_addr__h14584 ={32'd0, RTL__near_mem__dcache__cline_addr__h14583 }; 
  assign  RTL__near_mem__dcache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 = RTL__near_mem__dcache__dmem_not_imem &&! RTL__near_mem__dcache__soc_map$m_is_mem_addr || RTL__near_mem__dcache__rg_op ||! RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]||! RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL__near_mem__dcache__fabric_addr__h17243 ={32'd0, RTL__near_mem__dcache__rg_pa }; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [10:3]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [18:11]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [18:3]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [26:19]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [34:19]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [34:27]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [34:3]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [42:35]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [50:35]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [50:43]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [58:51]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:35]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:51]; 
  assign  RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 = RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:59]; 
  assign  RTL__near_mem__dcache__mem_req_wr_addr_awaddr__h2473 ={32'd0, RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [95:64]}; 
  assign  RTL__near_mem__dcache__pa_ctag__h4952 ={2'd0, RTL__near_mem__dcache__rg_addr [31:12]}; 
  assign  RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 = RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [21:0]== RTL__near_mem__dcache__pa_ctag__h4952 ; 
  assign  RTL__near_mem__dcache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 = RTL__near_mem__dcache__req_f3 [1:0]==2'b0|| RTL__near_mem__dcache__req_f3 [1:0]==2'b01&&! RTL__near_mem__dcache__req_addr [0]|| RTL__near_mem__dcache__req_f3 [1:0]==2'b10&& RTL__near_mem__dcache__req_addr [1:0]==2'b0|| RTL__near_mem__dcache__req_f3 [1:0]==2'b11&& RTL__near_mem__dcache__req_addr [2:0]==3'b0; 
  assign  RTL__near_mem__dcache__result__h11657 ={{56{ RTL__near_mem__dcache__word64094_BITS_15_TO_8__q18 [7]}}, RTL__near_mem__dcache__word64094_BITS_15_TO_8__q18 }; 
  assign  RTL__near_mem__dcache__result__h11685 ={{56{ RTL__near_mem__dcache__word64094_BITS_23_TO_16__q19 [7]}}, RTL__near_mem__dcache__word64094_BITS_23_TO_16__q19 }; 
  assign  RTL__near_mem__dcache__result__h11713 ={{56{ RTL__near_mem__dcache__word64094_BITS_31_TO_24__q21 [7]}}, RTL__near_mem__dcache__word64094_BITS_31_TO_24__q21 }; 
  assign  RTL__near_mem__dcache__result__h11741 ={{56{ RTL__near_mem__dcache__word64094_BITS_39_TO_32__q22 [7]}}, RTL__near_mem__dcache__word64094_BITS_39_TO_32__q22 }; 
  assign  RTL__near_mem__dcache__result__h11769 ={{56{ RTL__near_mem__dcache__word64094_BITS_47_TO_40__q25 [7]}}, RTL__near_mem__dcache__word64094_BITS_47_TO_40__q25 }; 
  assign  RTL__near_mem__dcache__result__h11797 ={{56{ RTL__near_mem__dcache__word64094_BITS_55_TO_48__q26 [7]}}, RTL__near_mem__dcache__word64094_BITS_55_TO_48__q26 }; 
  assign  RTL__near_mem__dcache__result__h11825 ={{56{ RTL__near_mem__dcache__word64094_BITS_63_TO_56__q28 [7]}}, RTL__near_mem__dcache__word64094_BITS_63_TO_56__q28 }; 
  assign  RTL__near_mem__dcache__result__h11870 ={56'd0, RTL__near_mem__dcache__word64__h5094 [7:0]}; 
  assign  RTL__near_mem__dcache__result__h11898 ={56'd0, RTL__near_mem__dcache__word64__h5094 [15:8]}; 
  assign  RTL__near_mem__dcache__result__h11926 ={56'd0, RTL__near_mem__dcache__word64__h5094 [23:16]}; 
  assign  RTL__near_mem__dcache__result__h11954 ={56'd0, RTL__near_mem__dcache__word64__h5094 [31:24]}; 
  assign  RTL__near_mem__dcache__result__h11982 ={56'd0, RTL__near_mem__dcache__word64__h5094 [39:32]}; 
  assign  RTL__near_mem__dcache__result__h12010 ={56'd0, RTL__near_mem__dcache__word64__h5094 [47:40]}; 
  assign  RTL__near_mem__dcache__result__h12038 ={56'd0, RTL__near_mem__dcache__word64__h5094 [55:48]}; 
  assign  RTL__near_mem__dcache__result__h12066 ={56'd0, RTL__near_mem__dcache__word64__h5094 [63:56]}; 
  assign  RTL__near_mem__dcache__result__h12111 ={{48{ RTL__near_mem__dcache__word64094_BITS_15_TO_0__q16 [15]}}, RTL__near_mem__dcache__word64094_BITS_15_TO_0__q16 }; 
  assign  RTL__near_mem__dcache__result__h12139 ={{48{ RTL__near_mem__dcache__word64094_BITS_31_TO_16__q20 [15]}}, RTL__near_mem__dcache__word64094_BITS_31_TO_16__q20 }; 
  assign  RTL__near_mem__dcache__result__h12167 ={{48{ RTL__near_mem__dcache__word64094_BITS_47_TO_32__q23 [15]}}, RTL__near_mem__dcache__word64094_BITS_47_TO_32__q23 }; 
  assign  RTL__near_mem__dcache__result__h12195 ={{48{ RTL__near_mem__dcache__word64094_BITS_63_TO_48__q27 [15]}}, RTL__near_mem__dcache__word64094_BITS_63_TO_48__q27 }; 
  assign  RTL__near_mem__dcache__result__h12236 ={48'd0, RTL__near_mem__dcache__word64__h5094 [15:0]}; 
  assign  RTL__near_mem__dcache__result__h12264 ={48'd0, RTL__near_mem__dcache__word64__h5094 [31:16]}; 
  assign  RTL__near_mem__dcache__result__h12292 ={48'd0, RTL__near_mem__dcache__word64__h5094 [47:32]}; 
  assign  RTL__near_mem__dcache__result__h12320 ={48'd0, RTL__near_mem__dcache__word64__h5094 [63:48]}; 
  assign  RTL__near_mem__dcache__result__h12361 ={{32{ RTL__near_mem__dcache__word64094_BITS_31_TO_0__q17 [31]}}, RTL__near_mem__dcache__word64094_BITS_31_TO_0__q17 }; 
  assign  RTL__near_mem__dcache__result__h12389 ={{32{ RTL__near_mem__dcache__word64094_BITS_63_TO_32__q24 [31]}}, RTL__near_mem__dcache__word64094_BITS_63_TO_32__q24 }; 
  assign  RTL__near_mem__dcache__result__h12428 ={32'd0, RTL__near_mem__dcache__word64__h5094 [31:0]}; 
  assign  RTL__near_mem__dcache__result__h12456 ={32'd0, RTL__near_mem__dcache__word64__h5094 [63:32]}; 
  assign  RTL__near_mem__dcache__result__h17654 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 }; 
  assign  RTL__near_mem__dcache__result__h17684 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 }; 
  assign  RTL__near_mem__dcache__result__h17711 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 }; 
  assign  RTL__near_mem__dcache__result__h17738 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 }; 
  assign  RTL__near_mem__dcache__result__h17765 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 }; 
  assign  RTL__near_mem__dcache__result__h17792 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 }; 
  assign  RTL__near_mem__dcache__result__h17819 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 }; 
  assign  RTL__near_mem__dcache__result__h17846 ={{56{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 [7]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 }; 
  assign  RTL__near_mem__dcache__result__h17890 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [10:3]}; 
  assign  RTL__near_mem__dcache__result__h17917 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [18:11]}; 
  assign  RTL__near_mem__dcache__result__h17944 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [26:19]}; 
  assign  RTL__near_mem__dcache__result__h17971 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [34:27]}; 
  assign  RTL__near_mem__dcache__result__h17998 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [42:35]}; 
  assign  RTL__near_mem__dcache__result__h18025 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [50:43]}; 
  assign  RTL__near_mem__dcache__result__h18052 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [58:51]}; 
  assign  RTL__near_mem__dcache__result__h18079 ={56'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:59]}; 
  assign  RTL__near_mem__dcache__result__h18123 ={{48{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 [15]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 }; 
  assign  RTL__near_mem__dcache__result__h18150 ={{48{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 [15]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 }; 
  assign  RTL__near_mem__dcache__result__h18177 ={{48{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 [15]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 }; 
  assign  RTL__near_mem__dcache__result__h18204 ={{48{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 [15]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 }; 
  assign  RTL__near_mem__dcache__result__h18244 ={48'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [18:3]}; 
  assign  RTL__near_mem__dcache__result__h18271 ={48'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [34:19]}; 
  assign  RTL__near_mem__dcache__result__h18298 ={48'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [50:35]}; 
  assign  RTL__near_mem__dcache__result__h18325 ={48'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:51]}; 
  assign  RTL__near_mem__dcache__result__h18365 ={{32{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 [31]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 }; 
  assign  RTL__near_mem__dcache__result__h18392 ={{32{ RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 [31]}}, RTL__near_mem__dcache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 }; 
  assign  RTL__near_mem__dcache__result__h18430 ={32'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [34:3]}; 
  assign  RTL__near_mem__dcache__result__h18457 ={32'd0, RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:35]}; 
  assign  RTL__near_mem__dcache__result__h5301 ={{56{ RTL__near_mem__dcache__word64094_BITS_7_TO_0__q15 [7]}}, RTL__near_mem__dcache__word64094_BITS_7_TO_0__q15 }; 
  assign  RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 = RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL__near_mem__dcache__shift_bits__h2487 ={ RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [66:64],3'b0}; 
  assign  RTL__near_mem__dcache__strobe64__h2637 =8'b00000001<< RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL__near_mem__dcache__strobe64__h2639 =8'b00000011<< RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL__near_mem__dcache__strobe64__h2641 =8'b00001111<< RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL__near_mem__dcache__word64094_BITS_15_TO_0__q16 = RTL__near_mem__dcache__word64__h5094 [15:0]; 
  assign  RTL__near_mem__dcache__word64094_BITS_15_TO_8__q18 = RTL__near_mem__dcache__word64__h5094 [15:8]; 
  assign  RTL__near_mem__dcache__word64094_BITS_23_TO_16__q19 = RTL__near_mem__dcache__word64__h5094 [23:16]; 
  assign  RTL__near_mem__dcache__word64094_BITS_31_TO_0__q17 = RTL__near_mem__dcache__word64__h5094 [31:0]; 
  assign  RTL__near_mem__dcache__word64094_BITS_31_TO_16__q20 = RTL__near_mem__dcache__word64__h5094 [31:16]; 
  assign  RTL__near_mem__dcache__word64094_BITS_31_TO_24__q21 = RTL__near_mem__dcache__word64__h5094 [31:24]; 
  assign  RTL__near_mem__dcache__word64094_BITS_39_TO_32__q22 = RTL__near_mem__dcache__word64__h5094 [39:32]; 
  assign  RTL__near_mem__dcache__word64094_BITS_47_TO_32__q23 = RTL__near_mem__dcache__word64__h5094 [47:32]; 
  assign  RTL__near_mem__dcache__word64094_BITS_47_TO_40__q25 = RTL__near_mem__dcache__word64__h5094 [47:40]; 
  assign  RTL__near_mem__dcache__word64094_BITS_55_TO_48__q26 = RTL__near_mem__dcache__word64__h5094 [55:48]; 
  assign  RTL__near_mem__dcache__word64094_BITS_63_TO_32__q24 = RTL__near_mem__dcache__word64__h5094 [63:32]; 
  assign  RTL__near_mem__dcache__word64094_BITS_63_TO_48__q27 = RTL__near_mem__dcache__word64__h5094 [63:48]; 
  assign  RTL__near_mem__dcache__word64094_BITS_63_TO_56__q28 = RTL__near_mem__dcache__word64__h5094 [63:56]; 
  assign  RTL__near_mem__dcache__word64094_BITS_7_TO_0__q15 = RTL__near_mem__dcache__word64__h5094 [7:0]; 
  assign  RTL__near_mem__dcache__word64__h5094 = RTL__near_mem__dcache__ram_word64_set$DOB & RTL__near_mem__dcache__y__h5337 ; 
  assign  RTL__near_mem__dcache__y__h5337 ={64{ RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 }}; 
  always @(  RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT  )
         begin 
             case ( RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL__near_mem__dcache__x__h2520  =3'b0;
              2 'b01: 
                  RTL__near_mem__dcache__x__h2520  =3'b001;
              2 'b10: 
                  RTL__near_mem__dcache__x__h2520  =3'b010;
              2 'b11: 
                  RTL__near_mem__dcache__x__h2520  =3'b011;endcase
         end
  always @(  RTL__near_mem__dcache__rg_f3  )
         begin 
             case ( RTL__near_mem__dcache__rg_f3 [1:0])
              2 'b0: 
                  RTL__near_mem__dcache__value__h17372  =3'b0;
              2 'b01: 
                  RTL__near_mem__dcache__value__h17372  =3'b001;
              2 'b10: 
                  RTL__near_mem__dcache__value__h17372  =3'b010;
              2 'd3: 
                  RTL__near_mem__dcache__value__h17372  =3'b011;endcase
         end
  always @(     RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT                or   RTL__near_mem__dcache__strobe64__h2637            or   RTL__near_mem__dcache__strobe64__h2639           or   RTL__near_mem__dcache__strobe64__h2641  )
         begin 
             case ( RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700  = RTL__near_mem__dcache__strobe64__h2637 ;
              2 'b01: 
                  RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700  = RTL__near_mem__dcache__strobe64__h2639 ;
              2 'b10: 
                  RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700  = RTL__near_mem__dcache__strobe64__h2641 ;
              2 'b11: 
                  RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700  =8'b11111111;endcase
         end
  always @(   RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT            or   RTL__near_mem__dcache___theResult___snd_fst__h2707  )
         begin 
             case ( RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [97:96])
              2 'b0,2'b01,2'b10: 
                  RTL__near_mem__dcache__mem_req_wr_data_wdata__h2699  = RTL__near_mem__dcache___theResult___snd_fst__h2707 ;
              2 'd3: 
                  RTL__near_mem__dcache__mem_req_wr_data_wdata__h2699  = RTL__near_mem__dcache__f_fabric_write_reqs$D_OUT [63:0];endcase
         end
  always @(      RTL__near_mem__dcache__rg_addr                  or   RTL__near_mem__dcache__result__h12111             or   RTL__near_mem__dcache__result__h12139            or   RTL__near_mem__dcache__result__h12167           or   RTL__near_mem__dcache__result__h12195  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__dcache__result__h12111 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__dcache__result__h12139 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__dcache__result__h12167 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__dcache__result__h12195 ;
              default : 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  =64'd0;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__ram_word64_set$DOB           or   RTL__near_mem__dcache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:16], RTL__near_mem__dcache__rg_st_amo_val [15:0]};
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:32], RTL__near_mem__dcache__rg_st_amo_val [15:0], RTL__near_mem__dcache__ram_word64_set$DOB [15:0]};
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:48], RTL__near_mem__dcache__rg_st_amo_val [15:0], RTL__near_mem__dcache__ram_word64_set$DOB [31:0]};
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__dcache__rg_st_amo_val [15:0], RTL__near_mem__dcache__ram_word64_set$DOB [47:0]};
              default : 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  = RTL__near_mem__dcache__ram_word64_set$DOB ;endcase
         end
  always @(          RTL__near_mem__dcache__rg_addr                          or   RTL__near_mem__dcache__result__h5301                 or   RTL__near_mem__dcache__result__h11657                or   RTL__near_mem__dcache__result__h11685               or   RTL__near_mem__dcache__result__h11713              or   RTL__near_mem__dcache__result__h11741             or   RTL__near_mem__dcache__result__h11769            or   RTL__near_mem__dcache__result__h11797           or   RTL__near_mem__dcache__result__h11825  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h5301 ;
              3 'h1: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11657 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11685 ;
              3 'h3: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11713 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11741 ;
              3 'h5: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11769 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11797 ;
              3 'h7: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__dcache__result__h11825 ;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__ram_word64_set$DOB           or   RTL__near_mem__dcache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:8], RTL__near_mem__dcache__rg_st_amo_val [7:0]};
              3 'h1: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:16], RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [7:0]};
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:24], RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [15:0]};
              3 'h3: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:32], RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [23:0]};
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:40], RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [31:0]};
              3 'h5: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:48], RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [39:0]};
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:56], RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [47:0]};
              3 'h7: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__dcache__rg_st_amo_val [7:0], RTL__near_mem__dcache__ram_word64_set$DOB [55:0]};endcase
         end
  always @(      RTL__near_mem__dcache__rg_addr                  or   RTL__near_mem__dcache__result__h18244             or   RTL__near_mem__dcache__result__h18271            or   RTL__near_mem__dcache__result__h18298           or   RTL__near_mem__dcache__result__h18325  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__dcache__result__h18244 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__dcache__result__h18271 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__dcache__result__h18298 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__dcache__result__h18325 ;
              default : 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  =64'd0;endcase
         end
  always @(      RTL__near_mem__dcache__rg_addr                  or   RTL__near_mem__dcache__result__h12236             or   RTL__near_mem__dcache__result__h12264            or   RTL__near_mem__dcache__result__h12292           or   RTL__near_mem__dcache__result__h12320  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__dcache__result__h12236 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__dcache__result__h12264 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__dcache__result__h12292 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__dcache__result__h12320 ;
              default : 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  =64'd0;endcase
         end
  always @(      RTL__near_mem__dcache__rg_addr                  or   RTL__near_mem__dcache__result__h18123             or   RTL__near_mem__dcache__result__h18150            or   RTL__near_mem__dcache__result__h18177           or   RTL__near_mem__dcache__result__h18204  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__dcache__result__h18123 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__dcache__result__h18150 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__dcache__result__h18177 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__dcache__result__h18204 ;
              default : 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  =64'd0;endcase
         end
  always @(          RTL__near_mem__dcache__rg_addr                          or   RTL__near_mem__dcache__result__h17890                 or   RTL__near_mem__dcache__result__h17917                or   RTL__near_mem__dcache__result__h17944               or   RTL__near_mem__dcache__result__h17971              or   RTL__near_mem__dcache__result__h17998             or   RTL__near_mem__dcache__result__h18025            or   RTL__near_mem__dcache__result__h18052           or   RTL__near_mem__dcache__result__h18079  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h17890 ;
              3 'h1: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h17917 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h17944 ;
              3 'h3: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h17971 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h17998 ;
              3 'h5: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h18025 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h18052 ;
              3 'h7: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__dcache__result__h18079 ;endcase
         end
  always @(          RTL__near_mem__dcache__rg_addr                          or   RTL__near_mem__dcache__result__h11870                 or   RTL__near_mem__dcache__result__h11898                or   RTL__near_mem__dcache__result__h11926               or   RTL__near_mem__dcache__result__h11954              or   RTL__near_mem__dcache__result__h11982             or   RTL__near_mem__dcache__result__h12010            or   RTL__near_mem__dcache__result__h12038           or   RTL__near_mem__dcache__result__h12066  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h11870 ;
              3 'h1: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h11898 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h11926 ;
              3 'h3: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h11954 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h11982 ;
              3 'h5: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h12010 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h12038 ;
              3 'h7: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__dcache__result__h12066 ;endcase
         end
  always @(          RTL__near_mem__dcache__rg_addr                          or   RTL__near_mem__dcache__result__h17654                 or   RTL__near_mem__dcache__result__h17684                or   RTL__near_mem__dcache__result__h17711               or   RTL__near_mem__dcache__result__h17738              or   RTL__near_mem__dcache__result__h17765             or   RTL__near_mem__dcache__result__h17792            or   RTL__near_mem__dcache__result__h17819           or   RTL__near_mem__dcache__result__h17846  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17654 ;
              3 'h1: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17684 ;
              3 'h2: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17711 ;
              3 'h3: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17738 ;
              3 'h4: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17765 ;
              3 'h5: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17792 ;
              3 'h6: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17819 ;
              3 'h7: 
                  RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__dcache__result__h17846 ;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__result__h18365           or   RTL__near_mem__dcache__result__h18392  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL__near_mem__dcache__result__h18365 ;
              3 'h4: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL__near_mem__dcache__result__h18392 ;
              default : 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  =64'd0;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__result__h18430           or   RTL__near_mem__dcache__result__h18457  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL__near_mem__dcache__result__h18430 ;
              3 'h4: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL__near_mem__dcache__result__h18457 ;
              default : 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  =64'd0;endcase
         end
  always @(          RTL__near_mem__dcache__rg_f3                          or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411                 or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439                or   RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29               or   RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT             or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427            or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447           or   RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  )
         begin 
             case ( RTL__near_mem__dcache__rg_f3 )
              3 'b0: 
                  RTL__near_mem__dcache__ld_val__h17594  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 ;
              3 'b001: 
                  RTL__near_mem__dcache__ld_val__h17594  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 ;
              3 'b010: 
                  RTL__near_mem__dcache__ld_val__h17594  = RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 ;
              3 'b011: 
                  RTL__near_mem__dcache__ld_val__h17594  =( RTL__near_mem__dcache__rg_addr [2:0]==3'h0) ?  RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:3]:64'd0;
              3 'b100: 
                  RTL__near_mem__dcache__ld_val__h17594  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 ;
              3 'b101: 
                  RTL__near_mem__dcache__ld_val__h17594  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 ;
              3 'b110: 
                  RTL__near_mem__dcache__ld_val__h17594  = RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 ;
              3 'd7: 
                  RTL__near_mem__dcache__ld_val__h17594  =64'd0;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__ram_word64_set$DOB           or   RTL__near_mem__dcache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL__near_mem__dcache__ram_word64_set$DOB [63:32], RTL__near_mem__dcache__rg_st_amo_val [31:0]};
              3 'h4: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL__near_mem__dcache__rg_st_amo_val [31:0], RTL__near_mem__dcache__ram_word64_set$DOB [31:0]};
              default : 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  = RTL__near_mem__dcache__ram_word64_set$DOB ;endcase
         end
  always @(       RTL__near_mem__dcache__rg_f3                    or   RTL__near_mem__dcache__ram_word64_set$DOB              or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157             or   RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167            or   RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31           or   RTL__near_mem__dcache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__dcache__rg_f3 )
              3 'b0: 
                  RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 ;
              3 'b001: 
                  RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__dcache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 ;
              3 'b010: 
                  RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 ;
              3 'b011: 
                  RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__dcache__rg_st_amo_val ;
              default : 
                  RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__dcache__ram_word64_set$DOB ;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__result__h12361           or   RTL__near_mem__dcache__result__h12389  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL__near_mem__dcache__result__h12361 ;
              3 'h4: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL__near_mem__dcache__result__h12389 ;
              default : 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  =64'd0;endcase
         end
  always @(    RTL__near_mem__dcache__rg_addr              or   RTL__near_mem__dcache__result__h12428           or   RTL__near_mem__dcache__result__h12456  )
         begin 
             case ( RTL__near_mem__dcache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL__near_mem__dcache__result__h12428 ;
              3 'h4: 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL__near_mem__dcache__result__h12456 ;
              default : 
                  RTL__near_mem__dcache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  =64'd0;endcase
         end
  always @( posedge  RTL__near_mem__dcache__CLK )
         begin 
             if ( RTL__near_mem__dcache__RST_N ==1'b0)
                 begin  
                     RTL__near_mem__dcache__cfg_verbosity  <=4'd0; 
                     RTL__near_mem__dcache__ctr_wr_rsps_pending_crg  <=4'd0; 
                     RTL__near_mem__dcache__rg_cset_in_cache  <=7'd0; 
                     RTL__near_mem__dcache__rg_lower_word32_full  <=1'd0; 
                     RTL__near_mem__dcache__rg_state  <=4'd0;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__dcache__cfg_verbosity$EN ) 
                         RTL__near_mem__dcache__cfg_verbosity  <= RTL__near_mem__dcache__cfg_verbosity$D_IN ;
                     if ( RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$EN ) 
                         RTL__near_mem__dcache__ctr_wr_rsps_pending_crg  <= RTL__near_mem__dcache__ctr_wr_rsps_pending_crg$D_IN ;
                     if ( RTL__near_mem__dcache__rg_cset_in_cache$EN ) 
                         RTL__near_mem__dcache__rg_cset_in_cache  <= RTL__near_mem__dcache__rg_cset_in_cache$D_IN ;
                     if ( RTL__near_mem__dcache__rg_lower_word32_full$EN ) 
                         RTL__near_mem__dcache__rg_lower_word32_full  <= RTL__near_mem__dcache__rg_lower_word32_full$D_IN ;
                     if ( RTL__near_mem__dcache__rg_state$EN ) 
                         RTL__near_mem__dcache__rg_state  <= RTL__near_mem__dcache__rg_state$D_IN ;
                 end 
             if ( RTL__near_mem__dcache__rg_addr$EN ) 
                 RTL__near_mem__dcache__rg_addr  <= RTL__near_mem__dcache__rg_addr$D_IN ;
             if ( RTL__near_mem__dcache__rg_error_during_refill$EN ) 
                 RTL__near_mem__dcache__rg_error_during_refill  <= RTL__near_mem__dcache__rg_error_during_refill$D_IN ;
             if ( RTL__near_mem__dcache__rg_exc_code$EN ) 
                 RTL__near_mem__dcache__rg_exc_code  <= RTL__near_mem__dcache__rg_exc_code$D_IN ;
             if ( RTL__near_mem__dcache__rg_f3$EN ) 
                 RTL__near_mem__dcache__rg_f3  <= RTL__near_mem__dcache__rg_f3$D_IN ;
             if ( RTL__near_mem__dcache__rg_ld_val$EN ) 
                 RTL__near_mem__dcache__rg_ld_val  <= RTL__near_mem__dcache__rg_ld_val$D_IN ;
             if ( RTL__near_mem__dcache__rg_lower_word32$EN ) 
                 RTL__near_mem__dcache__rg_lower_word32  <= RTL__near_mem__dcache__rg_lower_word32$D_IN ;
             if ( RTL__near_mem__dcache__rg_op$EN ) 
                 RTL__near_mem__dcache__rg_op  <= RTL__near_mem__dcache__rg_op$D_IN ;
             if ( RTL__near_mem__dcache__rg_pa$EN ) 
                 RTL__near_mem__dcache__rg_pa  <= RTL__near_mem__dcache__rg_pa$D_IN ;
             if ( RTL__near_mem__dcache__rg_pte_pa$EN ) 
                 RTL__near_mem__dcache__rg_pte_pa  <= RTL__near_mem__dcache__rg_pte_pa$D_IN ;
             if ( RTL__near_mem__dcache__rg_st_amo_val$EN ) 
                 RTL__near_mem__dcache__rg_st_amo_val  <= RTL__near_mem__dcache__rg_st_amo_val$D_IN ;
             if ( RTL__near_mem__dcache__rg_word64_set_in_cache$EN ) 
                 RTL__near_mem__dcache__rg_word64_set_in_cache  <= RTL__near_mem__dcache__rg_word64_set_in_cache$D_IN ;
         end
  always @( negedge  RTL__near_mem__dcache__CLK )
         begin #0;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__ctr_wr_rsps_pending_crg ==4'd15)
                     begin  
                         RTL__near_mem__dcache__v__h2948  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h2942  = RTL__near_mem__dcache__v__h2948 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__ctr_wr_rsps_pending_crg ==4'd15)$display("%0d: ERROR: CreditCounter: overflow", RTL__near_mem__dcache__v__h2942 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__ctr_wr_rsps_pending_crg ==4'd15)$finish(32'd1);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Addr { ","awid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awaddr: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__mem_req_wr_addr_awaddr__h2473 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlen: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awsize: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__x__h2520 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awburst: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlock: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awcache: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awprot: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awqos: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awregion: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awuser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("                       ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Data { ","wdata: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__mem_req_wr_data_wdata__h2699 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wstrb: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__mem_req_wr_data_wstrb__h2700 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wlast: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("True");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wuser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127&& RTL__near_mem__dcache__cfg_verbosity !=4'd0&&! RTL__near_mem__dcache__f_reset_reqs$D_OUT )
                     begin  
                         RTL__near_mem__dcache__v__h3848  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h3842  = RTL__near_mem__dcache__v__h3848 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127&& RTL__near_mem__dcache__cfg_verbosity !=4'd0&&! RTL__near_mem__dcache__f_reset_reqs$D_OUT )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL__near_mem__dcache__v__h3842 ,"D_MMU_Cache",$signed(32'd128),$signed(32'd1));
                      else $display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL__near_mem__dcache__v__h3842 ,"I_MMU_Cache",$signed(32'd128),$signed(32'd1));
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__f_reset_reqs$D_OUT )
                     begin  
                         RTL__near_mem__dcache__v__h3949  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h3943  = RTL__near_mem__dcache__v__h3949 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_reset && RTL__near_mem__dcache__rg_cset_in_cache ==7'd127&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__f_reset_reqs$D_OUT )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_reset: Flushed", RTL__near_mem__dcache__v__h3943 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_reset: Flushed", RTL__near_mem__dcache__v__h3943 ,"I_MMU_Cache");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h4098  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h4092  = RTL__near_mem__dcache__v__h4098 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL__near_mem__dcache__v__h4092 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_addr );
                      else $display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL__near_mem__dcache__v__h4092 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_addr );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        eaddr = {CTag 0x%0h  CSet 0x%0h  Word64 0x%0h  Byte 0x%0h}", RTL__near_mem__dcache__pa_ctag__h4952 , RTL__near_mem__dcache__rg_addr [11:5], RTL__near_mem__dcache__rg_addr [4:3], RTL__near_mem__dcache__rg_addr [2:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x: (state, tag):", RTL__near_mem__dcache__rg_addr [11:5]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" (");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22])$write("CTAG_CLEAN");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22])$write("CTAG_EMPTY");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22])$write(", 0x%0x", RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [21:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22])$write(", --");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(")");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__dcache__rg_addr [11:5], RTL__near_mem__dcache__rg_addr [4:3]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" 0x%0x", RTL__near_mem__dcache__ram_word64_set$DOB );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    TLB result: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_Xlate_Result { ","outcome: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_XLATE_OK");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","pa: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__rg_addr );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","exc_code: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'hA," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__dcache__dmem_not_imem &&! RTL__near_mem__dcache__soc_map$m_is_mem_addr && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => IO_REQ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$display("        Write-Cache-Hit: pa 0x%0h word64 0x%0h", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_st_amo_val );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        New Word64_Set:");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__dcache__rg_addr [11:5], RTL__near_mem__dcache__rg_addr [4:3]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write(" 0x%0x", RTL__near_mem__dcache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op &&(! RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]||! RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Miss: pa 0x%0h word64 0x%0h", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_st_amo_val );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Hit/Miss: eaddr 0x%0h word64 0x%0h", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_st_amo_val );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__rg_op && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        => rl_write_response");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     begin  
                         RTL__near_mem__dcache__v__h12540  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h12534  = RTL__near_mem__dcache__v__h12540 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL__near_mem__dcache__v__h12534 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__word64__h5094 ,64'd0);
                      else $display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL__near_mem__dcache__v__h12534 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__word64__h5094 ,64'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&& RTL__near_mem__dcache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )$display("        Read-hit: addr 0x%0h word64 0x%0h", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__word64__h5094 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__dcache__dmem_not_imem || RTL__near_mem__dcache__soc_map$m_is_mem_addr )&&! RTL__near_mem__dcache__rg_op &&(! RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB [22]||! RTL__near_mem__dcache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Read Miss: -> CACHE_START_REFILL.");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h14531  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h14525  = RTL__near_mem__dcache__v__h14531 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_start_cache_refill: ", RTL__near_mem__dcache__v__h14525 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_cache_refill: ", RTL__near_mem__dcache__v__h14525 ,"I_MMU_Cache");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    To fabric: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__cline_fabric_addr__h14584 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd3);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'b011);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    Victim way %0d; => CACHE_REFILL",1'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     begin  
                         RTL__near_mem__dcache__v__h15336  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h15330  = RTL__near_mem__dcache__v__h15336 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop:", RTL__near_mem__dcache__v__h15330 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_cache_refill_rsps_loop:", RTL__near_mem__dcache__v__h15330 ,"I_MMU_Cache");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rdata: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rresp: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rlast: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 &&! RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","ruser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h",1'd0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h15578  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h15572  = RTL__near_mem__dcache__v__h15578 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL__near_mem__dcache__v__h15572 ,"D_MMU_Cache", RTL__near_mem__dcache__access_exc_code__h2256 );
                      else $display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL__near_mem__dcache__v__h15572 ,"I_MMU_Cache", RTL__near_mem__dcache__access_exc_code__h2256 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]==2'd3&&( RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__dcache__rg_error_during_refill )&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => MODULE_EXCEPTION_RSP");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]==2'd3&& RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0&&! RTL__near_mem__dcache__rg_error_during_refill && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => CACHE_REREQ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$display("        Updating Cache word64_set 0x%0h, word64_in_cline %0d) old => new", RTL__near_mem__dcache__rg_word64_set_in_cache , RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__dcache__rg_addr [11:5], RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL__near_mem__dcache__ram_word64_set$DOB );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__dcache__rg_addr [11:5], RTL__near_mem__dcache__rg_word64_set_in_cache [1:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_rereq && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL__near_mem__dcache__rg_addr [11:5], RTL__near_mem__dcache__rg_addr [11:3]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h17191  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h17185  = RTL__near_mem__dcache__v__h17191 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL__near_mem__dcache__v__h17185 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_f3 , RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_pa );
                      else $display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL__near_mem__dcache__v__h17185 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_f3 , RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_pa );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__fabric_addr__h17243 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__value__h17372 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h17485  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h17479  = RTL__near_mem__dcache__v__h17485 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL__near_mem__dcache__v__h17479 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_pa );
                      else $display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL__near_mem__dcache__v__h17479 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_pa );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rdata: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rresp: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rlast: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","ruser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h18585  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h18579  = RTL__near_mem__dcache__v__h18585 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__dcache__v__h18579 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__ld_val__h17594 );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__dcache__v__h18579 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__ld_val__h17594 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h18692  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h18686  = RTL__near_mem__dcache__v__h18692 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL__near_mem__dcache__v__h18686 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL__near_mem__dcache__v__h18686 ,"I_MMU_Cache");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h18797  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h18791  = RTL__near_mem__dcache__v__h18797 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__dcache__v__h18791 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_ld_val );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__dcache__v__h18791 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_ld_val );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h18877  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h18871  = RTL__near_mem__dcache__v__h18877 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL__near_mem__dcache__v__h18871 ,"D_MMU_Cache", RTL__near_mem__dcache__rg_f3 , RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_pa , RTL__near_mem__dcache__rg_st_amo_val );
                      else $display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL__near_mem__dcache__v__h18871 ,"I_MMU_Cache", RTL__near_mem__dcache__rg_f3 , RTL__near_mem__dcache__rg_addr , RTL__near_mem__dcache__rg_pa , RTL__near_mem__dcache__rg_st_amo_val );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_io_write_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => rl_ST_AMO_response");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h19505  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h19499  = RTL__near_mem__dcache__v__h19505 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL__near_mem__dcache__v__h19499 ,"D_MMU_Cache",$unsigned( RTL__near_mem__dcache__b__h14485 ));
                      else $write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL__near_mem__dcache__v__h19499 ,"I_MMU_Cache",$unsigned( RTL__near_mem__dcache__b__h14485 ));
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","bresp: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","buser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     begin  
                         RTL__near_mem__dcache__v__h19466  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h19460  = RTL__near_mem__dcache__v__h19466 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL__near_mem__dcache__v__h19460 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL__near_mem__dcache__v__h19460 ,"I_MMU_Cache");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("    ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","bresp: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","buser: ");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h",1'd0," }");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h3483  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h3477  = RTL__near_mem__dcache__v__h3483 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__WILL_FIRE_RL_rl_start_reset && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__dcache__dmem_not_imem )$display("%0d: %s.rl_start_reset", RTL__near_mem__dcache__v__h3477 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_reset", RTL__near_mem__dcache__v__h3477 ,"I_MMU_Cache");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__dcache__v__h19852  =$stime;#0;
                     end  
             RTL__near_mem__dcache__v__h19846  = RTL__near_mem__dcache__v__h19852 /32'd10;
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("%0d: %m.req: op:", RTL__near_mem__dcache__v__h19846 );
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__req_op )$write("CACHE_ST");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__dcache__req_op )$write("CACHE_LD");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" f3:%0d addr:0x%0h st_value:0x%0h", RTL__near_mem__dcache__req_f3 , RTL__near_mem__dcache__req_addr , RTL__near_mem__dcache__req_st_value ,"\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    priv:");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__req_priv ==2'b0)$write("U");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__req_priv ==2'b01)$write("S");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__req_priv ==2'b11)$write("M");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__dcache__req_priv !=2'b0&& RTL__near_mem__dcache__req_priv !=2'b01&& RTL__near_mem__dcache__req_priv !=2'b11)$write("RESERVED");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" sstatus_SUM:%0d mstatus_MXR:%0d satp:0x%0h", RTL__near_mem__dcache__req_sstatus_SUM , RTL__near_mem__dcache__req_mstatus_MXR , RTL__near_mem__dcache__req_satp ,"\n");
             if ( RTL__near_mem__dcache__RST_N !=1'b0)
                 if ( RTL__near_mem__dcache__EN_req && RTL__near_mem__dcache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 && RTL__near_mem__dcache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL__near_mem__dcache__req_addr [11:5], RTL__near_mem__dcache__req_addr [11:3]);
         end
  assign  RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL__near_mem__dcache__rg_addr ; 
  assign  RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL__near_mem__dcache__rg_pa ;
      
    wire RTL__near_mem__f_reset_rsps__RST;
    wire RTL__near_mem__f_reset_rsps__CLK;
    wire RTL__near_mem__f_reset_rsps__ENQ;
    wire RTL__near_mem__f_reset_rsps__CLR;
    wire RTL__near_mem__f_reset_rsps__DEQ;
    wire RTL__near_mem__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;

    parameter RTL__near_mem__f_reset_rsps__guarded =1; 
    reg RTL__near_mem__f_reset_rsps__empty_reg ; 
    reg RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__FULL_N = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__EMPTY_N = RTL__near_mem__f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__near_mem__f_reset_rsps__CLK )
         begin 
             if ( RTL__near_mem__f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__near_mem__f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__near_mem__f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__f_reset_rsps__CLR )
                         begin  
                             RTL__near_mem__f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__near_mem__f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__f_reset_rsps__ENQ &&! RTL__near_mem__f_reset_rsps__DEQ )
                             begin  
                                 RTL__near_mem__f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__near_mem__f_reset_rsps__full_reg  <=! RTL__near_mem__f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if (! RTL__near_mem__f_reset_rsps__ENQ && RTL__near_mem__f_reset_rsps__DEQ )
                                 begin  
                                     RTL__near_mem__f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__near_mem__f_reset_rsps__empty_reg  <=! RTL__near_mem__f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__f_reset_rsps__CLK )
         begin : RTL__near_mem__f_reset_rsps__error_checks 
           reg RTL__near_mem__f_reset_rsps__deqerror , RTL__near_mem__f_reset_rsps__enqerror ; 
             RTL__near_mem__f_reset_rsps__deqerror  =0; 
             RTL__near_mem__f_reset_rsps__enqerror  =0;
             if ( RTL__near_mem__f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__f_reset_rsps__empty_reg && RTL__near_mem__f_reset_rsps__DEQ )
                         begin  
                             RTL__near_mem__f_reset_rsps__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__f_reset_rsps__full_reg && RTL__near_mem__f_reset_rsps__ENQ &&(! RTL__near_mem__f_reset_rsps__DEQ || RTL__near_mem__f_reset_rsps__guarded ))
                         begin  
                             RTL__near_mem__f_reset_rsps__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__empty_reg ;
    assign RTL__near_mem__f_reset_rsps__RST = RTL__near_mem__RST_N;
    assign RTL__near_mem__f_reset_rsps__CLK = RTL__near_mem__CLK;
    assign RTL__near_mem__f_reset_rsps__ENQ = RTL__near_mem__f_reset_rsps$ENQ;
    assign RTL__near_mem__f_reset_rsps__CLR = RTL__near_mem__f_reset_rsps$CLR;
    assign RTL__near_mem__f_reset_rsps__DEQ = RTL__near_mem__f_reset_rsps$DEQ;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__f_reset_rsps$EMPTY_N = RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
      
    
    parameter RTL__near_mem__icache__dmem_not_imem =1'b0; reg[63:0] RTL__near_mem__icache__word64 ; 
    wire[63:0] RTL__near_mem__icache__mem_master_araddr , RTL__near_mem__icache__mem_master_awaddr , RTL__near_mem__icache__mem_master_wdata , RTL__near_mem__icache__st_amo_val ; 
    wire[31:0] RTL__near_mem__icache__addr ; 
    wire[7:0] RTL__near_mem__icache__mem_master_arlen , RTL__near_mem__icache__mem_master_awlen , RTL__near_mem__icache__mem_master_wstrb ; 
    wire[3:0] RTL__near_mem__icache__exc_code , RTL__near_mem__icache__mem_master_arcache , RTL__near_mem__icache__mem_master_arid , RTL__near_mem__icache__mem_master_arqos , RTL__near_mem__icache__mem_master_arregion , RTL__near_mem__icache__mem_master_awcache , RTL__near_mem__icache__mem_master_awid , RTL__near_mem__icache__mem_master_awqos , RTL__near_mem__icache__mem_master_awregion ; 
    wire[2:0] RTL__near_mem__icache__mem_master_arprot , RTL__near_mem__icache__mem_master_arsize , RTL__near_mem__icache__mem_master_awprot , RTL__near_mem__icache__mem_master_awsize ; 
    wire[1:0] RTL__near_mem__icache__mem_master_arburst , RTL__near_mem__icache__mem_master_awburst ; 
    wire RTL__near_mem__icache__RDY_server_flush_request_put , RTL__near_mem__icache__RDY_server_flush_response_get , RTL__near_mem__icache__RDY_server_reset_request_put , RTL__near_mem__icache__RDY_server_reset_response_get , RTL__near_mem__icache__RDY_set_verbosity , RTL__near_mem__icache__RDY_tlb_flush , RTL__near_mem__icache__exc , RTL__near_mem__icache__mem_master_arlock , RTL__near_mem__icache__mem_master_arvalid , RTL__near_mem__icache__mem_master_awlock , RTL__near_mem__icache__mem_master_awvalid , RTL__near_mem__icache__mem_master_bready , RTL__near_mem__icache__mem_master_rready , RTL__near_mem__icache__mem_master_wlast , RTL__near_mem__icache__mem_master_wvalid , RTL__near_mem__icache__valid ; 
    wire[3:0] RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port0__write_1 , RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port1__write_1 , RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port2__read , RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port3__read ; 
    wire RTL__near_mem__icache__ctr_wr_rsps_pending_crg$EN_port2__write , RTL__near_mem__icache__dw_valid$whas ; reg[3:0] RTL__near_mem__icache__cfg_verbosity ; 
    wire[3:0] RTL__near_mem__icache__cfg_verbosity$D_IN ; 
    wire RTL__near_mem__icache__cfg_verbosity$EN ; reg[3:0] RTL__near_mem__icache__ctr_wr_rsps_pending_crg ; 
    wire[3:0] RTL__near_mem__icache__ctr_wr_rsps_pending_crg$D_IN ; 
    wire RTL__near_mem__icache__ctr_wr_rsps_pending_crg$EN ; reg[31:0] RTL__near_mem__icache__rg_addr ; 
    wire[31:0] RTL__near_mem__icache__rg_addr$D_IN ; 
    wire RTL__near_mem__icache__rg_addr$EN ; reg[6:0] RTL__near_mem__icache__rg_cset_in_cache ; 
    wire[6:0] RTL__near_mem__icache__rg_cset_in_cache$D_IN ; 
    wire RTL__near_mem__icache__rg_cset_in_cache$EN ; 
    reg RTL__near_mem__icache__rg_error_during_refill ; 
    wire RTL__near_mem__icache__rg_error_during_refill$D_IN , RTL__near_mem__icache__rg_error_during_refill$EN ; reg[3:0] RTL__near_mem__icache__rg_exc_code ; reg[3:0] RTL__near_mem__icache__rg_exc_code$D_IN ; 
    wire RTL__near_mem__icache__rg_exc_code$EN ; reg[2:0] RTL__near_mem__icache__rg_f3 ; 
    wire[2:0] RTL__near_mem__icache__rg_f3$D_IN ; 
    wire RTL__near_mem__icache__rg_f3$EN ; reg[63:0] RTL__near_mem__icache__rg_ld_val ; 
    wire[63:0] RTL__near_mem__icache__rg_ld_val$D_IN ; 
    wire RTL__near_mem__icache__rg_ld_val$EN ; reg[31:0] RTL__near_mem__icache__rg_lower_word32 ; 
    wire[31:0] RTL__near_mem__icache__rg_lower_word32$D_IN ; 
    wire RTL__near_mem__icache__rg_lower_word32$EN ; 
    reg RTL__near_mem__icache__rg_lower_word32_full ; 
    wire RTL__near_mem__icache__rg_lower_word32_full$D_IN , RTL__near_mem__icache__rg_lower_word32_full$EN ; 
    reg RTL__near_mem__icache__rg_op ; 
    wire RTL__near_mem__icache__rg_op$D_IN , RTL__near_mem__icache__rg_op$EN ; reg[31:0] RTL__near_mem__icache__rg_pa ; 
    wire[31:0] RTL__near_mem__icache__rg_pa$D_IN ; 
    wire RTL__near_mem__icache__rg_pa$EN ; reg[31:0] RTL__near_mem__icache__rg_pte_pa ; 
    wire[31:0] RTL__near_mem__icache__rg_pte_pa$D_IN ; 
    wire RTL__near_mem__icache__rg_pte_pa$EN ; reg[63:0] RTL__near_mem__icache__rg_st_amo_val ; 
    wire[63:0] RTL__near_mem__icache__rg_st_amo_val$D_IN ; 
    wire RTL__near_mem__icache__rg_st_amo_val$EN ; reg[3:0] RTL__near_mem__icache__rg_state ; reg[3:0] RTL__near_mem__icache__rg_state$D_IN ; 
    wire RTL__near_mem__icache__rg_state$EN ; reg[8:0] RTL__near_mem__icache__rg_word64_set_in_cache ; 
    wire[8:0] RTL__near_mem__icache__rg_word64_set_in_cache$D_IN ; 
    wire RTL__near_mem__icache__rg_word64_set_in_cache$EN ; 
    wire[98:0] RTL__near_mem__icache__f_fabric_write_reqs$D_IN , RTL__near_mem__icache__f_fabric_write_reqs$D_OUT ; 
    wire RTL__near_mem__icache__f_fabric_write_reqs$CLR , RTL__near_mem__icache__f_fabric_write_reqs$DEQ , RTL__near_mem__icache__f_fabric_write_reqs$EMPTY_N , RTL__near_mem__icache__f_fabric_write_reqs$ENQ , RTL__near_mem__icache__f_fabric_write_reqs$FULL_N ; 
    wire RTL__near_mem__icache__f_reset_reqs$CLR , RTL__near_mem__icache__f_reset_reqs$DEQ , RTL__near_mem__icache__f_reset_reqs$D_IN , RTL__near_mem__icache__f_reset_reqs$D_OUT , RTL__near_mem__icache__f_reset_reqs$EMPTY_N , RTL__near_mem__icache__f_reset_reqs$ENQ , RTL__near_mem__icache__f_reset_reqs$FULL_N ; 
    wire RTL__near_mem__icache__f_reset_rsps$CLR , RTL__near_mem__icache__f_reset_rsps$DEQ , RTL__near_mem__icache__f_reset_rsps$D_IN , RTL__near_mem__icache__f_reset_rsps$D_OUT , RTL__near_mem__icache__f_reset_rsps$EMPTY_N , RTL__near_mem__icache__f_reset_rsps$ENQ , RTL__near_mem__icache__f_reset_rsps$FULL_N ; 
    wire[96:0] RTL__near_mem__icache__master_xactor_f_rd_addr$D_IN , RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT ; 
    wire RTL__near_mem__icache__master_xactor_f_rd_addr$CLR , RTL__near_mem__icache__master_xactor_f_rd_addr$DEQ , RTL__near_mem__icache__master_xactor_f_rd_addr$EMPTY_N , RTL__near_mem__icache__master_xactor_f_rd_addr$ENQ , RTL__near_mem__icache__master_xactor_f_rd_addr$FULL_N ; 
    wire[70:0] RTL__near_mem__icache__master_xactor_f_rd_data$D_IN , RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT ; 
    wire RTL__near_mem__icache__master_xactor_f_rd_data$CLR , RTL__near_mem__icache__master_xactor_f_rd_data$DEQ , RTL__near_mem__icache__master_xactor_f_rd_data$EMPTY_N , RTL__near_mem__icache__master_xactor_f_rd_data$ENQ , RTL__near_mem__icache__master_xactor_f_rd_data$FULL_N ; 
    wire[96:0] RTL__near_mem__icache__master_xactor_f_wr_addr$D_IN , RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_addr$CLR , RTL__near_mem__icache__master_xactor_f_wr_addr$DEQ , RTL__near_mem__icache__master_xactor_f_wr_addr$EMPTY_N , RTL__near_mem__icache__master_xactor_f_wr_addr$ENQ , RTL__near_mem__icache__master_xactor_f_wr_addr$FULL_N ; 
    wire[72:0] RTL__near_mem__icache__master_xactor_f_wr_data$D_IN , RTL__near_mem__icache__master_xactor_f_wr_data$D_OUT ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_data$CLR , RTL__near_mem__icache__master_xactor_f_wr_data$DEQ , RTL__near_mem__icache__master_xactor_f_wr_data$EMPTY_N , RTL__near_mem__icache__master_xactor_f_wr_data$ENQ , RTL__near_mem__icache__master_xactor_f_wr_data$FULL_N ; 
    wire[5:0] RTL__near_mem__icache__master_xactor_f_wr_resp$D_IN , RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_resp$CLR , RTL__near_mem__icache__master_xactor_f_wr_resp$DEQ , RTL__near_mem__icache__master_xactor_f_wr_resp$EMPTY_N , RTL__near_mem__icache__master_xactor_f_wr_resp$ENQ , RTL__near_mem__icache__master_xactor_f_wr_resp$FULL_N ; 
    wire[22:0] RTL__near_mem__icache__ram_state_and_ctag_cset$DIA , RTL__near_mem__icache__ram_state_and_ctag_cset$DIB , RTL__near_mem__icache__ram_state_and_ctag_cset$DOB ; 
    wire[6:0] RTL__near_mem__icache__ram_state_and_ctag_cset$ADDRA , RTL__near_mem__icache__ram_state_and_ctag_cset$ADDRB ; 
    wire RTL__near_mem__icache__ram_state_and_ctag_cset$ENA , RTL__near_mem__icache__ram_state_and_ctag_cset$ENB , RTL__near_mem__icache__ram_state_and_ctag_cset$WEA , RTL__near_mem__icache__ram_state_and_ctag_cset$WEB ; reg[63:0] RTL__near_mem__icache__ram_word64_set$DIB ; reg[8:0] RTL__near_mem__icache__ram_word64_set$ADDRB ; 
    wire[63:0] RTL__near_mem__icache__ram_word64_set$DIA , RTL__near_mem__icache__ram_word64_set$DOB ; 
    wire[8:0] RTL__near_mem__icache__ram_word64_set$ADDRA ; 
    wire RTL__near_mem__icache__ram_word64_set$ENA , RTL__near_mem__icache__ram_word64_set$ENB , RTL__near_mem__icache__ram_word64_set$WEA , RTL__near_mem__icache__ram_word64_set$WEB ; 
    wire[63:0] RTL__near_mem__icache__soc_map$m_is_IO_addr_addr , RTL__near_mem__icache__soc_map$m_is_mem_addr_addr , RTL__near_mem__icache__soc_map$m_is_near_mem_IO_addr_addr ; 
    wire RTL__near_mem__icache__soc_map$m_is_mem_addr ; 
    wire RTL__near_mem__icache__CAN_FIRE_RL_rl_ST_AMO_response , RTL__near_mem__icache__CAN_FIRE_RL_rl_cache_refill_rsps_loop , RTL__near_mem__icache__CAN_FIRE_RL_rl_discard_write_rsp , RTL__near_mem__icache__CAN_FIRE_RL_rl_drive_exception_rsp , RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req , RTL__near_mem__icache__CAN_FIRE_RL_rl_io_read_req , RTL__near_mem__icache__CAN_FIRE_RL_rl_io_read_rsp , RTL__near_mem__icache__CAN_FIRE_RL_rl_io_write_req , RTL__near_mem__icache__CAN_FIRE_RL_rl_maintain_io_read_rsp , RTL__near_mem__icache__CAN_FIRE_RL_rl_probe_and_immed_rsp , RTL__near_mem__icache__CAN_FIRE_RL_rl_rereq , RTL__near_mem__icache__CAN_FIRE_RL_rl_reset , RTL__near_mem__icache__CAN_FIRE_RL_rl_start_cache_refill , RTL__near_mem__icache__CAN_FIRE_RL_rl_start_reset , RTL__near_mem__icache__CAN_FIRE_mem_master_m_arready , RTL__near_mem__icache__CAN_FIRE_mem_master_m_awready , RTL__near_mem__icache__CAN_FIRE_mem_master_m_bvalid , RTL__near_mem__icache__CAN_FIRE_mem_master_m_rvalid , RTL__near_mem__icache__CAN_FIRE_mem_master_m_wready , RTL__near_mem__icache__CAN_FIRE_req , RTL__near_mem__icache__CAN_FIRE_server_flush_request_put , RTL__near_mem__icache__CAN_FIRE_server_flush_response_get , RTL__near_mem__icache__CAN_FIRE_server_reset_request_put , RTL__near_mem__icache__CAN_FIRE_server_reset_response_get , RTL__near_mem__icache__CAN_FIRE_set_verbosity , RTL__near_mem__icache__CAN_FIRE_tlb_flush , RTL__near_mem__icache__WILL_FIRE_RL_rl_ST_AMO_response , RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop , RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp , RTL__near_mem__icache__WILL_FIRE_RL_rl_drive_exception_rsp , RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req , RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req , RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp , RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req , RTL__near_mem__icache__WILL_FIRE_RL_rl_maintain_io_read_rsp , RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp , RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq , RTL__near_mem__icache__WILL_FIRE_RL_rl_reset , RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill , RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset , RTL__near_mem__icache__WILL_FIRE_mem_master_m_arready , RTL__near_mem__icache__WILL_FIRE_mem_master_m_awready , RTL__near_mem__icache__WILL_FIRE_mem_master_m_bvalid , RTL__near_mem__icache__WILL_FIRE_mem_master_m_rvalid , RTL__near_mem__icache__WILL_FIRE_mem_master_m_wready , RTL__near_mem__icache__WILL_FIRE_req , RTL__near_mem__icache__WILL_FIRE_server_flush_request_put , RTL__near_mem__icache__WILL_FIRE_server_flush_response_get , RTL__near_mem__icache__WILL_FIRE_server_reset_request_put , RTL__near_mem__icache__WILL_FIRE_server_reset_response_get , RTL__near_mem__icache__WILL_FIRE_set_verbosity , RTL__near_mem__icache__WILL_FIRE_tlb_flush ; reg[63:0] RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2 ; 
    wire[98:0] RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__VAL_1 , RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
    wire[96:0] RTL__near_mem__icache__MUX_master_xactor_f_rd_addr$enq_1__VAL_1 , RTL__near_mem__icache__MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
    wire[22:0] RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ; 
    wire[8:0] RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_2 , RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_4 ; 
    wire[6:0] RTL__near_mem__icache__MUX_rg_cset_in_cache$write_1__VAL_1 ; 
    wire[3:0] RTL__near_mem__icache__MUX_rg_exc_code$write_1__VAL_1 , RTL__near_mem__icache__MUX_rg_state$write_1__VAL_1 , RTL__near_mem__icache__MUX_rg_state$write_1__VAL_4 , RTL__near_mem__icache__MUX_rg_state$write_1__VAL_7 , RTL__near_mem__icache__MUX_rg_state$write_1__VAL_9 ; 
    wire RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_1 , RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_2 , RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_3 , RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__SEL_1 , RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 , RTL__near_mem__icache__MUX_ram_word64_set$a_put_1__SEL_1 , RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2 , RTL__near_mem__icache__MUX_rg_error_during_refill$write_1__SEL_1 , RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_1 , RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_2 , RTL__near_mem__icache__MUX_rg_state$write_1__SEL_10 , RTL__near_mem__icache__MUX_rg_state$write_1__SEL_2 , RTL__near_mem__icache__MUX_rg_state$write_1__SEL_3 , RTL__near_mem__icache__MUX_rg_state$write_1__SEL_7 , RTL__near_mem__icache__MUX_rg_state$write_1__SEL_9 ; reg[31:0] RTL__near_mem__icache__v__h2948 ; reg[31:0] RTL__near_mem__icache__v__h3848 ; reg[31:0] RTL__near_mem__icache__v__h3949 ; reg[31:0] RTL__near_mem__icache__v__h4098 ; reg[31:0] RTL__near_mem__icache__v__h12540 ; reg[31:0] RTL__near_mem__icache__v__h14531 ; reg[31:0] RTL__near_mem__icache__v__h15336 ; reg[31:0] RTL__near_mem__icache__v__h15578 ; reg[31:0] RTL__near_mem__icache__v__h17191 ; reg[31:0] RTL__near_mem__icache__v__h17485 ; reg[31:0] RTL__near_mem__icache__v__h18585 ; reg[31:0] RTL__near_mem__icache__v__h18692 ; reg[31:0] RTL__near_mem__icache__v__h18797 ; reg[31:0] RTL__near_mem__icache__v__h18877 ; reg[31:0] RTL__near_mem__icache__v__h19505 ; reg[31:0] RTL__near_mem__icache__v__h19466 ; reg[31:0] RTL__near_mem__icache__v__h3483 ; reg[31:0] RTL__near_mem__icache__v__h19852 ; reg[31:0] RTL__near_mem__icache__v__h2942 ; reg[31:0] RTL__near_mem__icache__v__h3477 ; reg[31:0] RTL__near_mem__icache__v__h3842 ; reg[31:0] RTL__near_mem__icache__v__h3943 ; reg[31:0] RTL__near_mem__icache__v__h4092 ; reg[31:0] RTL__near_mem__icache__v__h12534 ; reg[31:0] RTL__near_mem__icache__v__h14525 ; reg[31:0] RTL__near_mem__icache__v__h15330 ; reg[31:0] RTL__near_mem__icache__v__h15572 ; reg[31:0] RTL__near_mem__icache__v__h17185 ; reg[31:0] RTL__near_mem__icache__v__h17479 ; reg[31:0] RTL__near_mem__icache__v__h18579 ; reg[31:0] RTL__near_mem__icache__v__h18686 ; reg[31:0] RTL__near_mem__icache__v__h18791 ; reg[31:0] RTL__near_mem__icache__v__h18871 ; reg[31:0] RTL__near_mem__icache__v__h19460 ; reg[31:0] RTL__near_mem__icache__v__h19499 ; reg[31:0] RTL__near_mem__icache__v__h19846 ; reg[63:0] RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 , RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 , RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 , RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 , RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 , RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 , RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 , RTL__near_mem__icache__ld_val__h17594 , RTL__near_mem__icache__mem_req_wr_data_wdata__h2699 ; reg[7:0] RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700 ; reg[2:0] RTL__near_mem__icache__value__h17372 , RTL__near_mem__icache__x__h2520 ; 
    wire[63:0] RTL__near_mem__icache___theResult___snd_fst__h2707 , RTL__near_mem__icache__cline_fabric_addr__h14584 , RTL__near_mem__icache__fabric_addr__h17243 , RTL__near_mem__icache__mem_req_wr_addr_awaddr__h2473 , RTL__near_mem__icache__result__h11657 , RTL__near_mem__icache__result__h11685 , RTL__near_mem__icache__result__h11713 , RTL__near_mem__icache__result__h11741 , RTL__near_mem__icache__result__h11769 , RTL__near_mem__icache__result__h11797 , RTL__near_mem__icache__result__h11825 , RTL__near_mem__icache__result__h11870 , RTL__near_mem__icache__result__h11898 , RTL__near_mem__icache__result__h11926 , RTL__near_mem__icache__result__h11954 , RTL__near_mem__icache__result__h11982 , RTL__near_mem__icache__result__h12010 , RTL__near_mem__icache__result__h12038 , RTL__near_mem__icache__result__h12066 , RTL__near_mem__icache__result__h12111 , RTL__near_mem__icache__result__h12139 , RTL__near_mem__icache__result__h12167 , RTL__near_mem__icache__result__h12195 , RTL__near_mem__icache__result__h12236 , RTL__near_mem__icache__result__h12264 , RTL__near_mem__icache__result__h12292 , RTL__near_mem__icache__result__h12320 , RTL__near_mem__icache__result__h12361 , RTL__near_mem__icache__result__h12389 , RTL__near_mem__icache__result__h12428 , RTL__near_mem__icache__result__h12456 , RTL__near_mem__icache__result__h17654 , RTL__near_mem__icache__result__h17684 , RTL__near_mem__icache__result__h17711 , RTL__near_mem__icache__result__h17738 , RTL__near_mem__icache__result__h17765 , RTL__near_mem__icache__result__h17792 , RTL__near_mem__icache__result__h17819 , RTL__near_mem__icache__result__h17846 , RTL__near_mem__icache__result__h17890 , RTL__near_mem__icache__result__h17917 , RTL__near_mem__icache__result__h17944 , RTL__near_mem__icache__result__h17971 , RTL__near_mem__icache__result__h17998 , RTL__near_mem__icache__result__h18025 , RTL__near_mem__icache__result__h18052 , RTL__near_mem__icache__result__h18079 , RTL__near_mem__icache__result__h18123 , RTL__near_mem__icache__result__h18150 , RTL__near_mem__icache__result__h18177 , RTL__near_mem__icache__result__h18204 , RTL__near_mem__icache__result__h18244 , RTL__near_mem__icache__result__h18271 , RTL__near_mem__icache__result__h18298 , RTL__near_mem__icache__result__h18325 , RTL__near_mem__icache__result__h18365 , RTL__near_mem__icache__result__h18392 , RTL__near_mem__icache__result__h18430 , RTL__near_mem__icache__result__h18457 , RTL__near_mem__icache__result__h5301 , RTL__near_mem__icache__word64__h5094 , RTL__near_mem__icache__y__h5337 ; 
    wire[31:0] RTL__near_mem__icache__cline_addr__h14583 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 , RTL__near_mem__icache__word64094_BITS_31_TO_0__q17 , RTL__near_mem__icache__word64094_BITS_63_TO_32__q24 ; 
    wire[21:0] RTL__near_mem__icache__pa_ctag__h4952 ; 
    wire[15:0] RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 , RTL__near_mem__icache__word64094_BITS_15_TO_0__q16 , RTL__near_mem__icache__word64094_BITS_31_TO_16__q20 , RTL__near_mem__icache__word64094_BITS_47_TO_32__q23 , RTL__near_mem__icache__word64094_BITS_63_TO_48__q27 ; 
    wire[7:0] RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 , RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 , RTL__near_mem__icache__strobe64__h2637 , RTL__near_mem__icache__strobe64__h2639 , RTL__near_mem__icache__strobe64__h2641 , RTL__near_mem__icache__word64094_BITS_15_TO_8__q18 , RTL__near_mem__icache__word64094_BITS_23_TO_16__q19 , RTL__near_mem__icache__word64094_BITS_31_TO_24__q21 , RTL__near_mem__icache__word64094_BITS_39_TO_32__q22 , RTL__near_mem__icache__word64094_BITS_47_TO_40__q25 , RTL__near_mem__icache__word64094_BITS_55_TO_48__q26 , RTL__near_mem__icache__word64094_BITS_63_TO_56__q28 , RTL__near_mem__icache__word64094_BITS_7_TO_0__q15 ; 
    wire[5:0] RTL__near_mem__icache__shift_bits__h2487 ; 
    wire[3:0] RTL__near_mem__icache__access_exc_code__h2256 , RTL__near_mem__icache__b__h14485 ; 
    wire RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 , RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 , RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 , RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 , RTL__near_mem__icache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 , RTL__near_mem__icache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 , RTL__near_mem__icache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 , RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 , RTL__near_mem__icache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 , RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 ; 
  assign  RTL__near_mem__icache__RDY_set_verbosity =1'd1; 
  assign  RTL__near_mem__icache__CAN_FIRE_set_verbosity =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_set_verbosity = RTL__near_mem__icache__EN_set_verbosity ; 
  assign  RTL__near_mem__icache__RDY_server_reset_request_put = RTL__near_mem__icache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__icache__CAN_FIRE_server_reset_request_put = RTL__near_mem__icache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__icache__WILL_FIRE_server_reset_request_put = RTL__near_mem__icache__EN_server_reset_request_put ; 
  assign  RTL__near_mem__icache__RDY_server_reset_response_get =! RTL__near_mem__icache__f_reset_rsps$D_OUT && RTL__near_mem__icache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__icache__CAN_FIRE_server_reset_response_get =! RTL__near_mem__icache__f_reset_rsps$D_OUT && RTL__near_mem__icache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__icache__WILL_FIRE_server_reset_response_get = RTL__near_mem__icache__EN_server_reset_response_get ; 
  assign  RTL__near_mem__icache__CAN_FIRE_req =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_req = RTL__near_mem__icache__EN_req ; 
  assign  RTL__near_mem__icache__valid = RTL__near_mem__icache__dw_valid$whas ; 
  assign  RTL__near_mem__icache__addr = RTL__near_mem__icache__rg_addr ; 
  always @(       RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_1                    or   RTL__near_mem__icache__ld_val__h17594              or   RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_2             or   RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2            or   RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_3           or   RTL__near_mem__icache__rg_ld_val  )
         begin 
             case (1'b1) 
              RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_1  : 
                  RTL__near_mem__icache__word64  = RTL__near_mem__icache__ld_val__h17594 ; 
              RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_2  : 
                  RTL__near_mem__icache__word64  = RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2 ; 
              RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_3  : 
                  RTL__near_mem__icache__word64  = RTL__near_mem__icache__rg_ld_val ;
              default : 
                  RTL__near_mem__icache__word64  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL__near_mem__icache__st_amo_val = RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_2  ? 64'd0: RTL__near_mem__icache__rg_st_amo_val ; 
  assign  RTL__near_mem__icache__exc = RTL__near_mem__icache__rg_state ==4'd4; 
  assign  RTL__near_mem__icache__exc_code = RTL__near_mem__icache__rg_exc_code ; 
  assign  RTL__near_mem__icache__RDY_server_flush_request_put = RTL__near_mem__icache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__icache__CAN_FIRE_server_flush_request_put = RTL__near_mem__icache__f_reset_reqs$FULL_N ; 
  assign  RTL__near_mem__icache__WILL_FIRE_server_flush_request_put = RTL__near_mem__icache__EN_server_flush_request_put ; 
  assign  RTL__near_mem__icache__RDY_server_flush_response_get = RTL__near_mem__icache__f_reset_rsps$D_OUT && RTL__near_mem__icache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__icache__CAN_FIRE_server_flush_response_get = RTL__near_mem__icache__f_reset_rsps$D_OUT && RTL__near_mem__icache__f_reset_rsps$EMPTY_N ; 
  assign  RTL__near_mem__icache__WILL_FIRE_server_flush_response_get = RTL__near_mem__icache__EN_server_flush_response_get ; 
  assign  RTL__near_mem__icache__RDY_tlb_flush =1'd1; 
  assign  RTL__near_mem__icache__CAN_FIRE_tlb_flush =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_tlb_flush = RTL__near_mem__icache__EN_tlb_flush ; 
  assign  RTL__near_mem__icache__mem_master_awvalid = RTL__near_mem__icache__master_xactor_f_wr_addr$EMPTY_N ; 
  assign  RTL__near_mem__icache__mem_master_awid = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [96:93]; 
  assign  RTL__near_mem__icache__mem_master_awaddr = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [92:29]; 
  assign  RTL__near_mem__icache__mem_master_awlen = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [28:21]; 
  assign  RTL__near_mem__icache__mem_master_awsize = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [20:18]; 
  assign  RTL__near_mem__icache__mem_master_awburst = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [17:16]; 
  assign  RTL__near_mem__icache__mem_master_awlock = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [15]; 
  assign  RTL__near_mem__icache__mem_master_awcache = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [14:11]; 
  assign  RTL__near_mem__icache__mem_master_awprot = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [10:8]; 
  assign  RTL__near_mem__icache__mem_master_awqos = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [7:4]; 
  assign  RTL__near_mem__icache__mem_master_awregion = RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT [3:0]; 
  assign  RTL__near_mem__icache__CAN_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL__near_mem__icache__mem_master_wvalid = RTL__near_mem__icache__master_xactor_f_wr_data$EMPTY_N ; 
  assign  RTL__near_mem__icache__mem_master_wdata = RTL__near_mem__icache__master_xactor_f_wr_data$D_OUT [72:9]; 
  assign  RTL__near_mem__icache__mem_master_wstrb = RTL__near_mem__icache__master_xactor_f_wr_data$D_OUT [8:1]; 
  assign  RTL__near_mem__icache__mem_master_wlast = RTL__near_mem__icache__master_xactor_f_wr_data$D_OUT [0]; 
  assign  RTL__near_mem__icache__CAN_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL__near_mem__icache__CAN_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL__near_mem__icache__mem_master_bready = RTL__near_mem__icache__master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL__near_mem__icache__mem_master_arvalid = RTL__near_mem__icache__master_xactor_f_rd_addr$EMPTY_N ; 
  assign  RTL__near_mem__icache__mem_master_arid = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [96:93]; 
  assign  RTL__near_mem__icache__mem_master_araddr = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [92:29]; 
  assign  RTL__near_mem__icache__mem_master_arlen = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [28:21]; 
  assign  RTL__near_mem__icache__mem_master_arsize = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [20:18]; 
  assign  RTL__near_mem__icache__mem_master_arburst = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [17:16]; 
  assign  RTL__near_mem__icache__mem_master_arlock = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [15]; 
  assign  RTL__near_mem__icache__mem_master_arcache = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [14:11]; 
  assign  RTL__near_mem__icache__mem_master_arprot = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [10:8]; 
  assign  RTL__near_mem__icache__mem_master_arqos = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [7:4]; 
  assign  RTL__near_mem__icache__mem_master_arregion = RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT [3:0]; 
  assign  RTL__near_mem__icache__CAN_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL__near_mem__icache__CAN_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL__near_mem__icache__mem_master_rready = RTL__near_mem__icache__master_xactor_f_rd_data$FULL_N ;  
    
    parameter RTL__near_mem__icache__f_fabric_write_reqs__width =1; parameter RTL__near_mem__icache__f_fabric_write_reqs__guarded =1; 
    reg RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
    reg RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; reg[ RTL__near_mem__icache__f_fabric_write_reqs__width -1:0] RTL__near_mem__icache__f_fabric_write_reqs__data0_reg ; reg[ RTL__near_mem__icache__f_fabric_write_reqs__width -1:0] RTL__near_mem__icache__f_fabric_write_reqs__data1_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__FULL_N = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__EMPTY_N = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__D_OUT = RTL__near_mem__icache__f_fabric_write_reqs__data0_reg ; 
    wire RTL__near_mem__icache__f_fabric_write_reqs__d0di =( RTL__near_mem__icache__f_fabric_write_reqs__ENQ &&! RTL__near_mem__icache__f_fabric_write_reqs__empty_reg )||( RTL__near_mem__icache__f_fabric_write_reqs__ENQ && RTL__near_mem__icache__f_fabric_write_reqs__DEQ && RTL__near_mem__icache__f_fabric_write_reqs__full_reg ); 
    wire RTL__near_mem__icache__f_fabric_write_reqs__d0d1 = RTL__near_mem__icache__f_fabric_write_reqs__DEQ &&! RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
    wire RTL__near_mem__icache__f_fabric_write_reqs__d0h =((! RTL__near_mem__icache__f_fabric_write_reqs__DEQ )&&(! RTL__near_mem__icache__f_fabric_write_reqs__ENQ ))||(! RTL__near_mem__icache__f_fabric_write_reqs__DEQ && RTL__near_mem__icache__f_fabric_write_reqs__empty_reg )||(! RTL__near_mem__icache__f_fabric_write_reqs__ENQ && RTL__near_mem__icache__f_fabric_write_reqs__full_reg ); 
    wire RTL__near_mem__icache__f_fabric_write_reqs__d1di = RTL__near_mem__icache__f_fabric_write_reqs__ENQ & RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__f_fabric_write_reqs__CLK )
         begin 
             if ( RTL__near_mem__icache__f_fabric_write_reqs__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__f_fabric_write_reqs__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__f_fabric_write_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__f_fabric_write_reqs__CLR )
                         begin  
                             RTL__near_mem__icache__f_fabric_write_reqs__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__f_fabric_write_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__f_fabric_write_reqs__ENQ &&! RTL__near_mem__icache__f_fabric_write_reqs__DEQ )
                             begin  
                                 RTL__near_mem__icache__f_fabric_write_reqs__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__f_fabric_write_reqs__full_reg  <=! RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__f_fabric_write_reqs__DEQ &&! RTL__near_mem__icache__f_fabric_write_reqs__ENQ )
                                 begin  
                                     RTL__near_mem__icache__f_fabric_write_reqs__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__f_fabric_write_reqs__empty_reg  <=! RTL__near_mem__icache__f_fabric_write_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__f_fabric_write_reqs__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__f_fabric_write_reqs__data0_reg  <={ RTL__near_mem__icache__f_fabric_write_reqs__width { RTL__near_mem__icache__f_fabric_write_reqs__d0di }}& RTL__near_mem__icache__f_fabric_write_reqs__D_IN |{ RTL__near_mem__icache__f_fabric_write_reqs__width { RTL__near_mem__icache__f_fabric_write_reqs__d0d1 }}& RTL__near_mem__icache__f_fabric_write_reqs__data1_reg |{ RTL__near_mem__icache__f_fabric_write_reqs__width { RTL__near_mem__icache__f_fabric_write_reqs__d0h }}& RTL__near_mem__icache__f_fabric_write_reqs__data0_reg ; 
                 RTL__near_mem__icache__f_fabric_write_reqs__data1_reg  <= RTL__near_mem__icache__f_fabric_write_reqs__d1di  ?  RTL__near_mem__icache__f_fabric_write_reqs__D_IN : RTL__near_mem__icache__f_fabric_write_reqs__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__f_fabric_write_reqs__CLK )
         begin : RTL__near_mem__icache__f_fabric_write_reqs__error_checks 
           reg RTL__near_mem__icache__f_fabric_write_reqs__deqerror , RTL__near_mem__icache__f_fabric_write_reqs__enqerror ; 
             RTL__near_mem__icache__f_fabric_write_reqs__deqerror  =0; 
             RTL__near_mem__icache__f_fabric_write_reqs__enqerror  =0;
             if ( RTL__near_mem__icache__f_fabric_write_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__f_fabric_write_reqs__empty_reg && RTL__near_mem__icache__f_fabric_write_reqs__DEQ )
                         begin  
                             RTL__near_mem__icache__f_fabric_write_reqs__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__f_fabric_write_reqs__full_reg && RTL__near_mem__icache__f_fabric_write_reqs__ENQ &&(! RTL__near_mem__icache__f_fabric_write_reqs__DEQ || RTL__near_mem__icache__f_fabric_write_reqs__guarded ))
                         begin  
                             RTL__near_mem__icache__f_fabric_write_reqs__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__empty_reg ;
    parameter RTL__near_mem__icache__f_reset_reqs__width =1; parameter RTL__near_mem__icache__f_reset_reqs__guarded =1; 
    reg RTL__near_mem__icache__f_reset_reqs__full_reg ; 
    reg RTL__near_mem__icache__f_reset_reqs__empty_reg ; reg[ RTL__near_mem__icache__f_reset_reqs__width -1:0] RTL__near_mem__icache__f_reset_reqs__data0_reg ; reg[ RTL__near_mem__icache__f_reset_reqs__width -1:0] RTL__near_mem__icache__f_reset_reqs__data1_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__FULL_N = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__EMPTY_N = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__D_OUT = RTL__near_mem__icache__f_reset_reqs__data0_reg ; 
    wire RTL__near_mem__icache__f_reset_reqs__d0di =( RTL__near_mem__icache__f_reset_reqs__ENQ &&! RTL__near_mem__icache__f_reset_reqs__empty_reg )||( RTL__near_mem__icache__f_reset_reqs__ENQ && RTL__near_mem__icache__f_reset_reqs__DEQ && RTL__near_mem__icache__f_reset_reqs__full_reg ); 
    wire RTL__near_mem__icache__f_reset_reqs__d0d1 = RTL__near_mem__icache__f_reset_reqs__DEQ &&! RTL__near_mem__icache__f_reset_reqs__full_reg ; 
    wire RTL__near_mem__icache__f_reset_reqs__d0h =((! RTL__near_mem__icache__f_reset_reqs__DEQ )&&(! RTL__near_mem__icache__f_reset_reqs__ENQ ))||(! RTL__near_mem__icache__f_reset_reqs__DEQ && RTL__near_mem__icache__f_reset_reqs__empty_reg )||(! RTL__near_mem__icache__f_reset_reqs__ENQ && RTL__near_mem__icache__f_reset_reqs__full_reg ); 
    wire RTL__near_mem__icache__f_reset_reqs__d1di = RTL__near_mem__icache__f_reset_reqs__ENQ & RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__f_reset_reqs__CLK )
         begin 
             if ( RTL__near_mem__icache__f_reset_reqs__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__f_reset_reqs__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__f_reset_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__f_reset_reqs__CLR )
                         begin  
                             RTL__near_mem__icache__f_reset_reqs__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__f_reset_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__f_reset_reqs__ENQ &&! RTL__near_mem__icache__f_reset_reqs__DEQ )
                             begin  
                                 RTL__near_mem__icache__f_reset_reqs__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__f_reset_reqs__full_reg  <=! RTL__near_mem__icache__f_reset_reqs__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__f_reset_reqs__DEQ &&! RTL__near_mem__icache__f_reset_reqs__ENQ )
                                 begin  
                                     RTL__near_mem__icache__f_reset_reqs__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__f_reset_reqs__empty_reg  <=! RTL__near_mem__icache__f_reset_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__f_reset_reqs__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__f_reset_reqs__data0_reg  <={ RTL__near_mem__icache__f_reset_reqs__width { RTL__near_mem__icache__f_reset_reqs__d0di }}& RTL__near_mem__icache__f_reset_reqs__D_IN |{ RTL__near_mem__icache__f_reset_reqs__width { RTL__near_mem__icache__f_reset_reqs__d0d1 }}& RTL__near_mem__icache__f_reset_reqs__data1_reg |{ RTL__near_mem__icache__f_reset_reqs__width { RTL__near_mem__icache__f_reset_reqs__d0h }}& RTL__near_mem__icache__f_reset_reqs__data0_reg ; 
                 RTL__near_mem__icache__f_reset_reqs__data1_reg  <= RTL__near_mem__icache__f_reset_reqs__d1di  ?  RTL__near_mem__icache__f_reset_reqs__D_IN : RTL__near_mem__icache__f_reset_reqs__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__f_reset_reqs__CLK )
         begin : RTL__near_mem__icache__f_reset_reqs__error_checks 
           reg RTL__near_mem__icache__f_reset_reqs__deqerror , RTL__near_mem__icache__f_reset_reqs__enqerror ; 
             RTL__near_mem__icache__f_reset_reqs__deqerror  =0; 
             RTL__near_mem__icache__f_reset_reqs__enqerror  =0;
             if ( RTL__near_mem__icache__f_reset_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__f_reset_reqs__empty_reg && RTL__near_mem__icache__f_reset_reqs__DEQ )
                         begin  
                             RTL__near_mem__icache__f_reset_reqs__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__f_reset_reqs__full_reg && RTL__near_mem__icache__f_reset_reqs__ENQ &&(! RTL__near_mem__icache__f_reset_reqs__DEQ || RTL__near_mem__icache__f_reset_reqs__guarded ))
                         begin  
                             RTL__near_mem__icache__f_reset_reqs__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__empty_reg ;
    parameter RTL__near_mem__icache__f_reset_rsps__width =1; parameter RTL__near_mem__icache__f_reset_rsps__guarded =1; 
    reg RTL__near_mem__icache__f_reset_rsps__full_reg ; 
    reg RTL__near_mem__icache__f_reset_rsps__empty_reg ; reg[ RTL__near_mem__icache__f_reset_rsps__width -1:0] RTL__near_mem__icache__f_reset_rsps__data0_reg ; reg[ RTL__near_mem__icache__f_reset_rsps__width -1:0] RTL__near_mem__icache__f_reset_rsps__data1_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__FULL_N = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__EMPTY_N = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__D_OUT = RTL__near_mem__icache__f_reset_rsps__data0_reg ; 
    wire RTL__near_mem__icache__f_reset_rsps__d0di =( RTL__near_mem__icache__f_reset_rsps__ENQ &&! RTL__near_mem__icache__f_reset_rsps__empty_reg )||( RTL__near_mem__icache__f_reset_rsps__ENQ && RTL__near_mem__icache__f_reset_rsps__DEQ && RTL__near_mem__icache__f_reset_rsps__full_reg ); 
    wire RTL__near_mem__icache__f_reset_rsps__d0d1 = RTL__near_mem__icache__f_reset_rsps__DEQ &&! RTL__near_mem__icache__f_reset_rsps__full_reg ; 
    wire RTL__near_mem__icache__f_reset_rsps__d0h =((! RTL__near_mem__icache__f_reset_rsps__DEQ )&&(! RTL__near_mem__icache__f_reset_rsps__ENQ ))||(! RTL__near_mem__icache__f_reset_rsps__DEQ && RTL__near_mem__icache__f_reset_rsps__empty_reg )||(! RTL__near_mem__icache__f_reset_rsps__ENQ && RTL__near_mem__icache__f_reset_rsps__full_reg ); 
    wire RTL__near_mem__icache__f_reset_rsps__d1di = RTL__near_mem__icache__f_reset_rsps__ENQ & RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__f_reset_rsps__CLK )
         begin 
             if ( RTL__near_mem__icache__f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__f_reset_rsps__CLR )
                         begin  
                             RTL__near_mem__icache__f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__f_reset_rsps__ENQ &&! RTL__near_mem__icache__f_reset_rsps__DEQ )
                             begin  
                                 RTL__near_mem__icache__f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__f_reset_rsps__full_reg  <=! RTL__near_mem__icache__f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__f_reset_rsps__DEQ &&! RTL__near_mem__icache__f_reset_rsps__ENQ )
                                 begin  
                                     RTL__near_mem__icache__f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__f_reset_rsps__empty_reg  <=! RTL__near_mem__icache__f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__f_reset_rsps__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__f_reset_rsps__data0_reg  <={ RTL__near_mem__icache__f_reset_rsps__width { RTL__near_mem__icache__f_reset_rsps__d0di }}& RTL__near_mem__icache__f_reset_rsps__D_IN |{ RTL__near_mem__icache__f_reset_rsps__width { RTL__near_mem__icache__f_reset_rsps__d0d1 }}& RTL__near_mem__icache__f_reset_rsps__data1_reg |{ RTL__near_mem__icache__f_reset_rsps__width { RTL__near_mem__icache__f_reset_rsps__d0h }}& RTL__near_mem__icache__f_reset_rsps__data0_reg ; 
                 RTL__near_mem__icache__f_reset_rsps__data1_reg  <= RTL__near_mem__icache__f_reset_rsps__d1di  ?  RTL__near_mem__icache__f_reset_rsps__D_IN : RTL__near_mem__icache__f_reset_rsps__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__f_reset_rsps__CLK )
         begin : RTL__near_mem__icache__f_reset_rsps__error_checks 
           reg RTL__near_mem__icache__f_reset_rsps__deqerror , RTL__near_mem__icache__f_reset_rsps__enqerror ; 
             RTL__near_mem__icache__f_reset_rsps__deqerror  =0; 
             RTL__near_mem__icache__f_reset_rsps__enqerror  =0;
             if ( RTL__near_mem__icache__f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__f_reset_rsps__empty_reg && RTL__near_mem__icache__f_reset_rsps__DEQ )
                         begin  
                             RTL__near_mem__icache__f_reset_rsps__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__f_reset_rsps__full_reg && RTL__near_mem__icache__f_reset_rsps__ENQ &&(! RTL__near_mem__icache__f_reset_rsps__DEQ || RTL__near_mem__icache__f_reset_rsps__guarded ))
                         begin  
                             RTL__near_mem__icache__f_reset_rsps__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__full_reg ; 
  assign  RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__empty_reg ;
    parameter RTL__near_mem__icache__master_xactor_f_rd_addr__width =1; parameter RTL__near_mem__icache__master_xactor_f_rd_addr__guarded =1; 
    reg RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
    reg RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; reg[ RTL__near_mem__icache__master_xactor_f_rd_addr__width -1:0] RTL__near_mem__icache__master_xactor_f_rd_addr__data0_reg ; reg[ RTL__near_mem__icache__master_xactor_f_rd_addr__width -1:0] RTL__near_mem__icache__master_xactor_f_rd_addr__data1_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__FULL_N = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__EMPTY_N = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__D_OUT = RTL__near_mem__icache__master_xactor_f_rd_addr__data0_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__d0di =( RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ &&! RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg )||( RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ && RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ && RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__d0d1 = RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ &&! RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__d0h =((! RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ )&&(! RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ ))||(! RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ && RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg )||(! RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ && RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_rd_addr__d1di = RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ & RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__master_xactor_f_rd_addr__CLK )
         begin 
             if ( RTL__near_mem__icache__master_xactor_f_rd_addr__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__master_xactor_f_rd_addr__CLR )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ &&! RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ )
                             begin  
                                 RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg  <=! RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ &&! RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ )
                                 begin  
                                     RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg  <=! RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_rd_addr__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__master_xactor_f_rd_addr__data0_reg  <={ RTL__near_mem__icache__master_xactor_f_rd_addr__width { RTL__near_mem__icache__master_xactor_f_rd_addr__d0di }}& RTL__near_mem__icache__master_xactor_f_rd_addr__D_IN |{ RTL__near_mem__icache__master_xactor_f_rd_addr__width { RTL__near_mem__icache__master_xactor_f_rd_addr__d0d1 }}& RTL__near_mem__icache__master_xactor_f_rd_addr__data1_reg |{ RTL__near_mem__icache__master_xactor_f_rd_addr__width { RTL__near_mem__icache__master_xactor_f_rd_addr__d0h }}& RTL__near_mem__icache__master_xactor_f_rd_addr__data0_reg ; 
                 RTL__near_mem__icache__master_xactor_f_rd_addr__data1_reg  <= RTL__near_mem__icache__master_xactor_f_rd_addr__d1di  ?  RTL__near_mem__icache__master_xactor_f_rd_addr__D_IN : RTL__near_mem__icache__master_xactor_f_rd_addr__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_rd_addr__CLK )
         begin : RTL__near_mem__icache__master_xactor_f_rd_addr__error_checks 
           reg RTL__near_mem__icache__master_xactor_f_rd_addr__deqerror , RTL__near_mem__icache__master_xactor_f_rd_addr__enqerror ; 
             RTL__near_mem__icache__master_xactor_f_rd_addr__deqerror  =0; 
             RTL__near_mem__icache__master_xactor_f_rd_addr__enqerror  =0;
             if ( RTL__near_mem__icache__master_xactor_f_rd_addr__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg && RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_rd_addr__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg && RTL__near_mem__icache__master_xactor_f_rd_addr__ENQ &&(! RTL__near_mem__icache__master_xactor_f_rd_addr__DEQ || RTL__near_mem__icache__master_xactor_f_rd_addr__guarded ))
                         begin  
                             RTL__near_mem__icache__master_xactor_f_rd_addr__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__empty_reg ;
    parameter RTL__near_mem__icache__master_xactor_f_rd_data__width =1; parameter RTL__near_mem__icache__master_xactor_f_rd_data__guarded =1; 
    reg RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
    reg RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; reg[ RTL__near_mem__icache__master_xactor_f_rd_data__width -1:0] RTL__near_mem__icache__master_xactor_f_rd_data__data0_reg ; reg[ RTL__near_mem__icache__master_xactor_f_rd_data__width -1:0] RTL__near_mem__icache__master_xactor_f_rd_data__data1_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__FULL_N = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__EMPTY_N = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__D_OUT = RTL__near_mem__icache__master_xactor_f_rd_data__data0_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_rd_data__d0di =( RTL__near_mem__icache__master_xactor_f_rd_data__ENQ &&! RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg )||( RTL__near_mem__icache__master_xactor_f_rd_data__ENQ && RTL__near_mem__icache__master_xactor_f_rd_data__DEQ && RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_rd_data__d0d1 = RTL__near_mem__icache__master_xactor_f_rd_data__DEQ &&! RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_rd_data__d0h =((! RTL__near_mem__icache__master_xactor_f_rd_data__DEQ )&&(! RTL__near_mem__icache__master_xactor_f_rd_data__ENQ ))||(! RTL__near_mem__icache__master_xactor_f_rd_data__DEQ && RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg )||(! RTL__near_mem__icache__master_xactor_f_rd_data__ENQ && RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_rd_data__d1di = RTL__near_mem__icache__master_xactor_f_rd_data__ENQ & RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__master_xactor_f_rd_data__CLK )
         begin 
             if ( RTL__near_mem__icache__master_xactor_f_rd_data__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__master_xactor_f_rd_data__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__master_xactor_f_rd_data__CLR )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__master_xactor_f_rd_data__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__master_xactor_f_rd_data__ENQ &&! RTL__near_mem__icache__master_xactor_f_rd_data__DEQ )
                             begin  
                                 RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__master_xactor_f_rd_data__full_reg  <=! RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__master_xactor_f_rd_data__DEQ &&! RTL__near_mem__icache__master_xactor_f_rd_data__ENQ )
                                 begin  
                                     RTL__near_mem__icache__master_xactor_f_rd_data__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg  <=! RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_rd_data__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__master_xactor_f_rd_data__data0_reg  <={ RTL__near_mem__icache__master_xactor_f_rd_data__width { RTL__near_mem__icache__master_xactor_f_rd_data__d0di }}& RTL__near_mem__icache__master_xactor_f_rd_data__D_IN |{ RTL__near_mem__icache__master_xactor_f_rd_data__width { RTL__near_mem__icache__master_xactor_f_rd_data__d0d1 }}& RTL__near_mem__icache__master_xactor_f_rd_data__data1_reg |{ RTL__near_mem__icache__master_xactor_f_rd_data__width { RTL__near_mem__icache__master_xactor_f_rd_data__d0h }}& RTL__near_mem__icache__master_xactor_f_rd_data__data0_reg ; 
                 RTL__near_mem__icache__master_xactor_f_rd_data__data1_reg  <= RTL__near_mem__icache__master_xactor_f_rd_data__d1di  ?  RTL__near_mem__icache__master_xactor_f_rd_data__D_IN : RTL__near_mem__icache__master_xactor_f_rd_data__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_rd_data__CLK )
         begin : RTL__near_mem__icache__master_xactor_f_rd_data__error_checks 
           reg RTL__near_mem__icache__master_xactor_f_rd_data__deqerror , RTL__near_mem__icache__master_xactor_f_rd_data__enqerror ; 
             RTL__near_mem__icache__master_xactor_f_rd_data__deqerror  =0; 
             RTL__near_mem__icache__master_xactor_f_rd_data__enqerror  =0;
             if ( RTL__near_mem__icache__master_xactor_f_rd_data__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg && RTL__near_mem__icache__master_xactor_f_rd_data__DEQ )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_rd_data__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__master_xactor_f_rd_data__full_reg && RTL__near_mem__icache__master_xactor_f_rd_data__ENQ &&(! RTL__near_mem__icache__master_xactor_f_rd_data__DEQ || RTL__near_mem__icache__master_xactor_f_rd_data__guarded ))
                         begin  
                             RTL__near_mem__icache__master_xactor_f_rd_data__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__empty_reg ;
    parameter RTL__near_mem__icache__master_xactor_f_wr_addr__width =1; parameter RTL__near_mem__icache__master_xactor_f_wr_addr__guarded =1; 
    reg RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
    reg RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; reg[ RTL__near_mem__icache__master_xactor_f_wr_addr__width -1:0] RTL__near_mem__icache__master_xactor_f_wr_addr__data0_reg ; reg[ RTL__near_mem__icache__master_xactor_f_wr_addr__width -1:0] RTL__near_mem__icache__master_xactor_f_wr_addr__data1_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__FULL_N = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__EMPTY_N = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__D_OUT = RTL__near_mem__icache__master_xactor_f_wr_addr__data0_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__d0di =( RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ &&! RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg )||( RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ && RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ && RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__d0d1 = RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ &&! RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__d0h =((! RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ )&&(! RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ ))||(! RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ && RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg )||(! RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ && RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_wr_addr__d1di = RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ & RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_addr__CLK )
         begin 
             if ( RTL__near_mem__icache__master_xactor_f_wr_addr__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__master_xactor_f_wr_addr__CLR )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ &&! RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ )
                             begin  
                                 RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg  <=! RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ &&! RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ )
                                 begin  
                                     RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg  <=! RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_addr__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__master_xactor_f_wr_addr__data0_reg  <={ RTL__near_mem__icache__master_xactor_f_wr_addr__width { RTL__near_mem__icache__master_xactor_f_wr_addr__d0di }}& RTL__near_mem__icache__master_xactor_f_wr_addr__D_IN |{ RTL__near_mem__icache__master_xactor_f_wr_addr__width { RTL__near_mem__icache__master_xactor_f_wr_addr__d0d1 }}& RTL__near_mem__icache__master_xactor_f_wr_addr__data1_reg |{ RTL__near_mem__icache__master_xactor_f_wr_addr__width { RTL__near_mem__icache__master_xactor_f_wr_addr__d0h }}& RTL__near_mem__icache__master_xactor_f_wr_addr__data0_reg ; 
                 RTL__near_mem__icache__master_xactor_f_wr_addr__data1_reg  <= RTL__near_mem__icache__master_xactor_f_wr_addr__d1di  ?  RTL__near_mem__icache__master_xactor_f_wr_addr__D_IN : RTL__near_mem__icache__master_xactor_f_wr_addr__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_addr__CLK )
         begin : RTL__near_mem__icache__master_xactor_f_wr_addr__error_checks 
           reg RTL__near_mem__icache__master_xactor_f_wr_addr__deqerror , RTL__near_mem__icache__master_xactor_f_wr_addr__enqerror ; 
             RTL__near_mem__icache__master_xactor_f_wr_addr__deqerror  =0; 
             RTL__near_mem__icache__master_xactor_f_wr_addr__enqerror  =0;
             if ( RTL__near_mem__icache__master_xactor_f_wr_addr__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg && RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_addr__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg && RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ &&(! RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ || RTL__near_mem__icache__master_xactor_f_wr_addr__guarded ))
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_addr__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__empty_reg ;
    parameter RTL__near_mem__icache__master_xactor_f_wr_data__width =1; parameter RTL__near_mem__icache__master_xactor_f_wr_data__guarded =1; 
    reg RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
    reg RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; reg[ RTL__near_mem__icache__master_xactor_f_wr_data__width -1:0] RTL__near_mem__icache__master_xactor_f_wr_data__data0_reg ; reg[ RTL__near_mem__icache__master_xactor_f_wr_data__width -1:0] RTL__near_mem__icache__master_xactor_f_wr_data__data1_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__FULL_N = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__EMPTY_N = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__D_OUT = RTL__near_mem__icache__master_xactor_f_wr_data__data0_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_data__d0di =( RTL__near_mem__icache__master_xactor_f_wr_data__ENQ &&! RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg )||( RTL__near_mem__icache__master_xactor_f_wr_data__ENQ && RTL__near_mem__icache__master_xactor_f_wr_data__DEQ && RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_wr_data__d0d1 = RTL__near_mem__icache__master_xactor_f_wr_data__DEQ &&! RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_data__d0h =((! RTL__near_mem__icache__master_xactor_f_wr_data__DEQ )&&(! RTL__near_mem__icache__master_xactor_f_wr_data__ENQ ))||(! RTL__near_mem__icache__master_xactor_f_wr_data__DEQ && RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg )||(! RTL__near_mem__icache__master_xactor_f_wr_data__ENQ && RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_wr_data__d1di = RTL__near_mem__icache__master_xactor_f_wr_data__ENQ & RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_data__CLK )
         begin 
             if ( RTL__near_mem__icache__master_xactor_f_wr_data__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__master_xactor_f_wr_data__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__master_xactor_f_wr_data__CLR )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__master_xactor_f_wr_data__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__master_xactor_f_wr_data__ENQ &&! RTL__near_mem__icache__master_xactor_f_wr_data__DEQ )
                             begin  
                                 RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__master_xactor_f_wr_data__full_reg  <=! RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__master_xactor_f_wr_data__DEQ &&! RTL__near_mem__icache__master_xactor_f_wr_data__ENQ )
                                 begin  
                                     RTL__near_mem__icache__master_xactor_f_wr_data__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg  <=! RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_data__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__master_xactor_f_wr_data__data0_reg  <={ RTL__near_mem__icache__master_xactor_f_wr_data__width { RTL__near_mem__icache__master_xactor_f_wr_data__d0di }}& RTL__near_mem__icache__master_xactor_f_wr_data__D_IN |{ RTL__near_mem__icache__master_xactor_f_wr_data__width { RTL__near_mem__icache__master_xactor_f_wr_data__d0d1 }}& RTL__near_mem__icache__master_xactor_f_wr_data__data1_reg |{ RTL__near_mem__icache__master_xactor_f_wr_data__width { RTL__near_mem__icache__master_xactor_f_wr_data__d0h }}& RTL__near_mem__icache__master_xactor_f_wr_data__data0_reg ; 
                 RTL__near_mem__icache__master_xactor_f_wr_data__data1_reg  <= RTL__near_mem__icache__master_xactor_f_wr_data__d1di  ?  RTL__near_mem__icache__master_xactor_f_wr_data__D_IN : RTL__near_mem__icache__master_xactor_f_wr_data__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_data__CLK )
         begin : RTL__near_mem__icache__master_xactor_f_wr_data__error_checks 
           reg RTL__near_mem__icache__master_xactor_f_wr_data__deqerror , RTL__near_mem__icache__master_xactor_f_wr_data__enqerror ; 
             RTL__near_mem__icache__master_xactor_f_wr_data__deqerror  =0; 
             RTL__near_mem__icache__master_xactor_f_wr_data__enqerror  =0;
             if ( RTL__near_mem__icache__master_xactor_f_wr_data__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg && RTL__near_mem__icache__master_xactor_f_wr_data__DEQ )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_data__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__master_xactor_f_wr_data__full_reg && RTL__near_mem__icache__master_xactor_f_wr_data__ENQ &&(! RTL__near_mem__icache__master_xactor_f_wr_data__DEQ || RTL__near_mem__icache__master_xactor_f_wr_data__guarded ))
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_data__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__empty_reg ;
    parameter RTL__near_mem__icache__master_xactor_f_wr_resp__width =1; parameter RTL__near_mem__icache__master_xactor_f_wr_resp__guarded =1; 
    reg RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
    reg RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; reg[ RTL__near_mem__icache__master_xactor_f_wr_resp__width -1:0] RTL__near_mem__icache__master_xactor_f_wr_resp__data0_reg ; reg[ RTL__near_mem__icache__master_xactor_f_wr_resp__width -1:0] RTL__near_mem__icache__master_xactor_f_wr_resp__data1_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__FULL_N = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__EMPTY_N = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__D_OUT = RTL__near_mem__icache__master_xactor_f_wr_resp__data0_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__d0di =( RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ &&! RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg )||( RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ && RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ && RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__d0d1 = RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ &&! RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__d0h =((! RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ )&&(! RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ ))||(! RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ && RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg )||(! RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ && RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ); 
    wire RTL__near_mem__icache__master_xactor_f_wr_resp__d1di = RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ & RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_resp__CLK )
         begin 
             if ( RTL__near_mem__icache__master_xactor_f_wr_resp__RST ==1'b0)
                 begin  
                     RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg  <=1'b0; 
                     RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__master_xactor_f_wr_resp__CLR )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg  <=1'b0; 
                             RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ &&! RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ )
                             begin  
                                 RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg  <=1'b1; 
                                 RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg  <=! RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ;
                             end 
                          else 
                             if ( RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ &&! RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ )
                                 begin  
                                     RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg  <=1'b1; 
                                     RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg  <=! RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_resp__CLK )
         begin 
             begin  
                 RTL__near_mem__icache__master_xactor_f_wr_resp__data0_reg  <={ RTL__near_mem__icache__master_xactor_f_wr_resp__width { RTL__near_mem__icache__master_xactor_f_wr_resp__d0di }}& RTL__near_mem__icache__master_xactor_f_wr_resp__D_IN |{ RTL__near_mem__icache__master_xactor_f_wr_resp__width { RTL__near_mem__icache__master_xactor_f_wr_resp__d0d1 }}& RTL__near_mem__icache__master_xactor_f_wr_resp__data1_reg |{ RTL__near_mem__icache__master_xactor_f_wr_resp__width { RTL__near_mem__icache__master_xactor_f_wr_resp__d0h }}& RTL__near_mem__icache__master_xactor_f_wr_resp__data0_reg ; 
                 RTL__near_mem__icache__master_xactor_f_wr_resp__data1_reg  <= RTL__near_mem__icache__master_xactor_f_wr_resp__d1di  ?  RTL__near_mem__icache__master_xactor_f_wr_resp__D_IN : RTL__near_mem__icache__master_xactor_f_wr_resp__data1_reg ;
             end 
         end
  always @( posedge  RTL__near_mem__icache__master_xactor_f_wr_resp__CLK )
         begin : RTL__near_mem__icache__master_xactor_f_wr_resp__error_checks 
           reg RTL__near_mem__icache__master_xactor_f_wr_resp__deqerror , RTL__near_mem__icache__master_xactor_f_wr_resp__enqerror ; 
             RTL__near_mem__icache__master_xactor_f_wr_resp__deqerror  =0; 
             RTL__near_mem__icache__master_xactor_f_wr_resp__enqerror  =0;
             if ( RTL__near_mem__icache__master_xactor_f_wr_resp__RST ==!1'b0)
                 begin 
                     if (! RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg && RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ )
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_resp__deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg && RTL__near_mem__icache__master_xactor_f_wr_resp__ENQ &&(! RTL__near_mem__icache__master_xactor_f_wr_resp__DEQ || RTL__near_mem__icache__master_xactor_f_wr_resp__guarded ))
                         begin  
                             RTL__near_mem__icache__master_xactor_f_wr_resp__enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__full_reg ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__empty_reg ;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__f_fabric_write_reqs$D_IN = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_fabric_write_reqs$ENQ = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_fabric_write_reqs$DEQ = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__f_fabric_write_reqs$EMPTY_N = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$D_IN = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$ENQ = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$DEQ = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$CLR = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$D_OUT = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$FULL_N = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_reqs$EMPTY_N = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__f_reset_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__f_reset_rsps$ENQ = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__f_reset_rsps$DEQ = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__dcache__f_reset_rsps$CLR = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_rsps$D_OUT = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_rsps$FULL_N = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__f_reset_rsps$EMPTY_N = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__f_reset_rsps__RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__f_reset_rsps__CLK = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__f_reset_rsps__RST = RTL__near_mem__dcache__RST_N;
    assign RTL__near_mem__dcache__f_reset_rsps__D_IN = RTL__near_mem__dcache__f_reset_rsps$D_IN;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr__ENQ = RTL__near_mem__dcache__master_xactor_f_rd_addr$ENQ;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr__DEQ = RTL__near_mem__dcache__master_xactor_f_rd_addr$DEQ;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr__CLR = RTL__near_mem__dcache__master_xactor_f_rd_addr$CLR;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr$FULL_N = RTL__near_mem__dcache__master_xactor_f_rd_addr__FULL_N;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr$EMPTY_N = RTL__near_mem__dcache__master_xactor_f_rd_addr__EMPTY_N;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr$D_OUT = RTL__near_mem__dcache__master_xactor_f_rd_addr__D_OUT;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_rd_addr$EMPTY_N = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_rd_data$D_IN = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_rd_data$CLR = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_rd_data$D_OUT = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_rd_data$FULL_N = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_rd_data$EMPTY_N = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_addr$ENQ = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_addr$DEQ = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_addr$D_OUT = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_addr$FULL_N = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_addr$EMPTY_N = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data$D_IN = RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data__CLK = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data__RST = RTL__near_mem__dcache__RST_N;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data__D_IN = RTL__near_mem__dcache__master_xactor_f_wr_data$D_IN;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data__ENQ = RTL__near_mem__dcache__master_xactor_f_wr_data$ENQ;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data__DEQ = RTL__near_mem__dcache__master_xactor_f_wr_data$DEQ;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data__CLR = RTL__near_mem__dcache__master_xactor_f_wr_data$CLR;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data$FULL_N = RTL__near_mem__dcache__master_xactor_f_wr_data__FULL_N;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data$EMPTY_N = RTL__near_mem__dcache__master_xactor_f_wr_data__EMPTY_N;
    assign RTL__near_mem__dcache__master_xactor_f_wr_data$D_OUT = RTL__near_mem__dcache__master_xactor_f_wr_data__D_OUT;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$D_IN = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$ENQ = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$DEQ = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$CLR = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$D_OUT = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$FULL_N = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache__master_xactor_f_wr_resp$EMPTY_N = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$D_IN = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$ENQ = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$DEQ = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$CLR = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$D_OUT = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$FULL_N = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__icache__f_fabric_write_reqs$EMPTY_N = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__f_fabric_write_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache__f_reset_reqs$D_IN = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__f_reset_reqs$ENQ = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__f_reset_reqs$CLR = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__f_reset_reqs$D_OUT = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__f_reset_reqs$EMPTY_N = RTL__near_mem__icache__f_reset_reqs__RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache__f_reset_reqs__CLK = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__f_reset_reqs__RST = RTL__near_mem__icache__RST_N;
    assign RTL__near_mem__icache__f_reset_reqs__D_IN = RTL__near_mem__icache__f_reset_reqs$D_IN;
    assign RTL__near_mem__icache__f_reset_reqs__ENQ = RTL__near_mem__icache__f_reset_reqs$ENQ;
    assign RTL__near_mem__icache__f_reset_rsps__DEQ = RTL__near_mem__icache__f_reset_rsps$DEQ;
    assign RTL__near_mem__icache__f_reset_rsps__CLR = RTL__near_mem__icache__f_reset_rsps$CLR;
    assign RTL__near_mem__icache__f_reset_rsps$FULL_N = RTL__near_mem__icache__f_reset_rsps__FULL_N;
    assign RTL__near_mem__icache__f_reset_rsps$EMPTY_N = RTL__near_mem__icache__f_reset_rsps__EMPTY_N;
    assign RTL__near_mem__icache__f_reset_rsps$D_OUT = RTL__near_mem__icache__f_reset_rsps__D_OUT;
    assign RTL__near_mem__icache__f_reset_rsps$CLR = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__f_reset_rsps$D_OUT = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__icache__f_reset_rsps$FULL_N = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__f_reset_rsps__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$D_IN = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$ENQ = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$DEQ = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$CLR = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$D_OUT = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$FULL_N = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_addr$EMPTY_N = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_addr__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_data$D_IN = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_data$DEQ = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_data$CLR = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_data$FULL_N = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_rd_data$EMPTY_N = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_rd_data__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr__CLK = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr__RST = RTL__near_mem__icache__RST_N;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr__D_IN = RTL__near_mem__icache__master_xactor_f_wr_addr$D_IN;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr__ENQ = RTL__near_mem__icache__master_xactor_f_wr_addr$ENQ;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr__DEQ = RTL__near_mem__icache__master_xactor_f_wr_addr$DEQ;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr__CLR = RTL__near_mem__icache__master_xactor_f_wr_addr$CLR;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr$FULL_N = RTL__near_mem__icache__master_xactor_f_wr_addr__FULL_N;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr$EMPTY_N = RTL__near_mem__icache__master_xactor_f_wr_addr__EMPTY_N;
    assign RTL__near_mem__icache__master_xactor_f_wr_addr$D_OUT = RTL__near_mem__icache__master_xactor_f_wr_addr__D_OUT;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_addr__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_data$D_IN = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_data$ENQ = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_data$DEQ = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_data$CLR = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_data$D_OUT = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_data$EMPTY_N = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_data__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_resp$ENQ = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_resp$DEQ = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_resp$CLR = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_resp$FULL_N = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__icache__master_xactor_f_wr_resp$EMPTY_N = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__master_xactor_f_wr_resp__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
      
    
    reg[ RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R ; reg[ RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R ; reg[ RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R2 ; reg[ RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R2 ; parameter RTL__near_mem__icache__ram_state_and_ctag_cset__PIPELINED =0; parameter RTL__near_mem__icache__ram_state_and_ctag_cset__ADDR_WIDTH =1; parameter RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH =1; parameter RTL__near_mem__icache__ram_state_and_ctag_cset__MEMSIZE =1; (* RTL__near_mem__icache__ram_state_and_ctag_cset__keep *)
    wire[ RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__arb1 ; (* RTL__near_mem__icache__ram_state_and_ctag_cset__keep *)
    wire[ RTL__near_mem__icache__ram_state_and_ctag_cset__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_state_and_ctag_cset__arb2 ; 
  always @( posedge  RTL__near_mem__icache__ram_state_and_ctag_cset__CLKA )
         begin 
             if ( RTL__near_mem__icache__ram_state_and_ctag_cset__ENA )
                 begin 
                     if ( RTL__near_mem__icache__ram_state_and_ctag_cset__WEA )
                         begin  
                             RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R  <= RTL__near_mem__icache__ram_state_and_ctag_cset__DIA ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R  <= RTL__near_mem__icache__ram_state_and_ctag_cset__arb1 ;
                         end 
                 end  
             RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R2  <= RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R ;
         end
  always @( posedge  RTL__near_mem__icache__ram_state_and_ctag_cset__CLKB )
         begin 
             if ( RTL__near_mem__icache__ram_state_and_ctag_cset__ENB )
                 begin 
                     if ( RTL__near_mem__icache__ram_state_and_ctag_cset__WEB )
                         begin  
                             RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R  <= RTL__near_mem__icache__ram_state_and_ctag_cset__DIB ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R  <= RTL__near_mem__icache__ram_state_and_ctag_cset__arb2 ;
                         end 
                 end  
             RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R2  <= RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R ;
         end
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset__DOA =( RTL__near_mem__icache__ram_state_and_ctag_cset__PIPELINED ) ?  RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R2 : RTL__near_mem__icache__ram_state_and_ctag_cset__DOA_R ; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset__DOB =( RTL__near_mem__icache__ram_state_and_ctag_cset__PIPELINED ) ?  RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R2 : RTL__near_mem__icache__ram_state_and_ctag_cset__DOB_R ;
    reg[ RTL__near_mem__icache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_word64_set__DOA_R ; reg[ RTL__near_mem__icache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_word64_set__DOB_R ; reg[ RTL__near_mem__icache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_word64_set__DOA_R2 ; reg[ RTL__near_mem__icache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_word64_set__DOB_R2 ; parameter RTL__near_mem__icache__ram_word64_set__PIPELINED =0; parameter RTL__near_mem__icache__ram_word64_set__ADDR_WIDTH =1; parameter RTL__near_mem__icache__ram_word64_set__DATA_WIDTH =1; parameter RTL__near_mem__icache__ram_word64_set__MEMSIZE =1; (* RTL__near_mem__icache__ram_word64_set__keep *)
    wire[ RTL__near_mem__icache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_word64_set__arb1 ; (* RTL__near_mem__icache__ram_word64_set__keep *)
    wire[ RTL__near_mem__icache__ram_word64_set__DATA_WIDTH -1:0] RTL__near_mem__icache__ram_word64_set__arb2 ; 
  always @( posedge  RTL__near_mem__icache__ram_word64_set__CLKA )
         begin 
             if ( RTL__near_mem__icache__ram_word64_set__ENA )
                 begin 
                     if ( RTL__near_mem__icache__ram_word64_set__WEA )
                         begin  
                             RTL__near_mem__icache__ram_word64_set__DOA_R  <= RTL__near_mem__icache__ram_word64_set__DIA ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__icache__ram_word64_set__DOA_R  <= RTL__near_mem__icache__ram_word64_set__arb1 ;
                         end 
                 end  
             RTL__near_mem__icache__ram_word64_set__DOA_R2  <= RTL__near_mem__icache__ram_word64_set__DOA_R ;
         end
  always @( posedge  RTL__near_mem__icache__ram_word64_set__CLKB )
         begin 
             if ( RTL__near_mem__icache__ram_word64_set__ENB )
                 begin 
                     if ( RTL__near_mem__icache__ram_word64_set__WEB )
                         begin  
                             RTL__near_mem__icache__ram_word64_set__DOB_R  <= RTL__near_mem__icache__ram_word64_set__DIB ;
                         end 
                      else 
                         begin  
                             RTL__near_mem__icache__ram_word64_set__DOB_R  <= RTL__near_mem__icache__ram_word64_set__arb2 ;
                         end 
                 end  
             RTL__near_mem__icache__ram_word64_set__DOB_R2  <= RTL__near_mem__icache__ram_word64_set__DOB_R ;
         end
  assign  RTL__near_mem__icache__ram_word64_set__DOA =( RTL__near_mem__icache__ram_word64_set__PIPELINED ) ?  RTL__near_mem__icache__ram_word64_set__DOA_R2 : RTL__near_mem__icache__ram_word64_set__DOA_R ; 
  assign  RTL__near_mem__icache__ram_word64_set__DOB =( RTL__near_mem__icache__ram_word64_set__PIPELINED ) ?  RTL__near_mem__icache__ram_word64_set__DOB_R2 : RTL__near_mem__icache__ram_word64_set__DOB_R ;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__CLKA = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__ENA = RTL__near_mem__dcache__ram_state_and_ctag_cset$ENA;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__WEA = RTL__near_mem__dcache__ram_state_and_ctag_cset$WEA;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDRA = RTL__near_mem__dcache__ram_state_and_ctag_cset$ADDRA;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__DIA = RTL__near_mem__dcache__ram_state_and_ctag_cset$DIA;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__CLKB = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__ENB = RTL__near_mem__dcache__ram_state_and_ctag_cset$ENB;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__WEB = RTL__near_mem__dcache__ram_state_and_ctag_cset$WEB;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__ADDRB = RTL__near_mem__dcache__ram_state_and_ctag_cset$ADDRB;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset__DIB = RTL__near_mem__dcache__ram_state_and_ctag_cset$DIB;
    assign RTL__near_mem__dcache__ram_state_and_ctag_cset$DOB = RTL__near_mem__dcache__ram_state_and_ctag_cset__DOB;
    assign RTL__near_mem__dcache__ram_word64_set__CLKA = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__ram_word64_set__ENA = RTL__near_mem__dcache__ram_word64_set$ENA;
    assign RTL__near_mem__dcache__ram_word64_set__WEA = RTL__near_mem__dcache__ram_word64_set$WEA;
    assign RTL__near_mem__dcache__ram_word64_set__ADDRA = RTL__near_mem__dcache__ram_word64_set$ADDRA;
    assign RTL__near_mem__dcache__ram_word64_set__DIA = RTL__near_mem__dcache__ram_word64_set$DIA;
    assign RTL__near_mem__dcache__ram_word64_set__CLKB = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__ram_word64_set__ENB = RTL__near_mem__dcache__ram_word64_set$ENB;
    assign RTL__near_mem__dcache__ram_word64_set__WEB = RTL__near_mem__dcache__ram_word64_set$WEB;
    assign RTL__near_mem__dcache__ram_word64_set__ADDRB = RTL__near_mem__dcache__ram_word64_set$ADDRB;
    assign RTL__near_mem__dcache__ram_word64_set__DIB = RTL__near_mem__dcache__ram_word64_set$DIB;
    assign RTL__near_mem__dcache__ram_word64_set$DOB = RTL__near_mem__dcache__ram_word64_set__DOB;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__CLKA = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__ENA = RTL__near_mem__icache__ram_state_and_ctag_cset$ENA;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__WEA = RTL__near_mem__icache__ram_state_and_ctag_cset$WEA;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__ADDRA = RTL__near_mem__icache__ram_state_and_ctag_cset$ADDRA;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__DIA = RTL__near_mem__icache__ram_state_and_ctag_cset$DIA;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__CLKB = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__ENB = RTL__near_mem__icache__ram_state_and_ctag_cset$ENB;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__WEB = RTL__near_mem__icache__ram_state_and_ctag_cset$WEB;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__ADDRB = RTL__near_mem__icache__ram_state_and_ctag_cset$ADDRB;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset__DIB = RTL__near_mem__icache__ram_state_and_ctag_cset$DIB;
    assign RTL__near_mem__icache__ram_state_and_ctag_cset$DOB = RTL__near_mem__icache__ram_state_and_ctag_cset__DOB;
    assign RTL__near_mem__icache__ram_word64_set__CLKA = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__ram_word64_set__ENA = RTL__near_mem__icache__ram_word64_set$ENA;
    assign RTL__near_mem__icache__ram_word64_set__WEA = RTL__near_mem__icache__ram_word64_set$WEA;
    assign RTL__near_mem__icache__ram_word64_set__ADDRA = RTL__near_mem__icache__ram_word64_set$ADDRA;
    assign RTL__near_mem__icache__ram_word64_set__DIA = RTL__near_mem__icache__ram_word64_set$DIA;
    assign RTL__near_mem__icache__ram_word64_set__CLKB = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__ram_word64_set__ENB = RTL__near_mem__icache__ram_word64_set$ENB;
    assign RTL__near_mem__icache__ram_word64_set__WEB = RTL__near_mem__icache__ram_word64_set$WEB;
    assign RTL__near_mem__icache__ram_word64_set__ADDRB = RTL__near_mem__icache__ram_word64_set$ADDRB;
    assign RTL__near_mem__icache__ram_word64_set__DIB = RTL__near_mem__icache__ram_word64_set$DIB;
    assign RTL__near_mem__icache__ram_word64_set$DOB = RTL__near_mem__icache__ram_word64_set__DOB;
      
    
    wire[63:0] RTL__near_mem__icache__soc_map__m_boot_rom_addr_base , RTL__near_mem__icache__soc_map__m_boot_rom_addr_lim , RTL__near_mem__icache__soc_map__m_boot_rom_addr_size , RTL__near_mem__icache__soc_map__m_mem0_controller_addr_base , RTL__near_mem__icache__soc_map__m_mem0_controller_addr_lim , RTL__near_mem__icache__soc_map__m_mem0_controller_addr_size , RTL__near_mem__icache__soc_map__m_mtvec_reset_value , RTL__near_mem__icache__soc_map__m_near_mem_io_addr_base , RTL__near_mem__icache__soc_map__m_near_mem_io_addr_lim , RTL__near_mem__icache__soc_map__m_near_mem_io_addr_size , RTL__near_mem__icache__soc_map__m_nmivec_reset_value , RTL__near_mem__icache__soc_map__m_pc_reset_value , RTL__near_mem__icache__soc_map__m_plic_addr_base , RTL__near_mem__icache__soc_map__m_plic_addr_lim , RTL__near_mem__icache__soc_map__m_plic_addr_size , RTL__near_mem__icache__soc_map__m_tcm_addr_base , RTL__near_mem__icache__soc_map__m_tcm_addr_lim , RTL__near_mem__icache__soc_map__m_tcm_addr_size , RTL__near_mem__icache__soc_map__m_uart0_addr_base , RTL__near_mem__icache__soc_map__m_uart0_addr_lim , RTL__near_mem__icache__soc_map__m_uart0_addr_size ; 
    wire RTL__near_mem__icache__soc_map__m_is_IO_addr , RTL__near_mem__icache__soc_map__m_is_mem_addr , RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr ; 
  assign  RTL__near_mem__icache__soc_map__m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL__near_mem__icache__soc_map__m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL__near_mem__icache__soc_map__m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL__near_mem__icache__soc_map__m_plic_addr_base =64'h000000000C000000; 
  assign  RTL__near_mem__icache__soc_map__m_plic_addr_size =64'h0000000000400000; 
  assign  RTL__near_mem__icache__soc_map__m_plic_addr_lim =64'd205520896; 
  assign  RTL__near_mem__icache__soc_map__m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL__near_mem__icache__soc_map__m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL__near_mem__icache__soc_map__m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL__near_mem__icache__soc_map__m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL__near_mem__icache__soc_map__m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL__near_mem__icache__soc_map__m_boot_rom_addr_lim =64'd8192; 
  assign  RTL__near_mem__icache__soc_map__m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL__near_mem__icache__soc_map__m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL__near_mem__icache__soc_map__m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL__near_mem__icache__soc_map__m_tcm_addr_base =64'h0; 
  assign  RTL__near_mem__icache__soc_map__m_tcm_addr_size =64'd0; 
  assign  RTL__near_mem__icache__soc_map__m_tcm_addr_lim =64'd0; 
  assign  RTL__near_mem__icache__soc_map__m_is_mem_addr = RTL__near_mem__icache__soc_map__m_is_mem_addr_addr >=64'h0000000000001000&& RTL__near_mem__icache__soc_map__m_is_mem_addr_addr <64'd8192|| RTL__near_mem__icache__soc_map__m_is_mem_addr_addr >=64'h0000000080000000&& RTL__near_mem__icache__soc_map__m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL__near_mem__icache__soc_map__m_is_IO_addr = RTL__near_mem__icache__soc_map__m_is_IO_addr_addr >=64'h0000000002000000&& RTL__near_mem__icache__soc_map__m_is_IO_addr_addr <64'd33603584|| RTL__near_mem__icache__soc_map__m_is_IO_addr_addr >=64'h000000000C000000&& RTL__near_mem__icache__soc_map__m_is_IO_addr_addr <64'd205520896|| RTL__near_mem__icache__soc_map__m_is_IO_addr_addr >=64'h00000000C0000000&& RTL__near_mem__icache__soc_map__m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr = RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL__near_mem__icache__soc_map__m_pc_reset_value =64'h0000000000001000; 
  assign  RTL__near_mem__icache__soc_map__m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL__near_mem__icache__soc_map__m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
     
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req = RTL__near_mem__icache__f_fabric_write_reqs$EMPTY_N && RTL__near_mem__icache__master_xactor_f_wr_addr$FULL_N && RTL__near_mem__icache__master_xactor_f_wr_data$FULL_N ; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req = RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_reset =( RTL__near_mem__icache__rg_cset_in_cache !=7'd127|| RTL__near_mem__icache__f_reset_reqs$EMPTY_N && RTL__near_mem__icache__f_reset_rsps$FULL_N )&& RTL__near_mem__icache__rg_state ==4'd1; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_reset = RTL__near_mem__icache__CAN_FIRE_RL_rl_reset ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_probe_and_immed_rsp =( RTL__near_mem__icache__dmem_not_imem &&! RTL__near_mem__icache__soc_map$m_is_mem_addr ||! RTL__near_mem__icache__rg_op || RTL__near_mem__icache__f_fabric_write_reqs$FULL_N )&& RTL__near_mem__icache__rg_state ==4'd3; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp = RTL__near_mem__icache__CAN_FIRE_RL_rl_probe_and_immed_rsp &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_start_cache_refill = RTL__near_mem__icache__master_xactor_f_rd_addr$FULL_N && RTL__near_mem__icache__rg_state ==4'd8&& RTL__near_mem__icache__b__h14485 ==4'd0; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill = RTL__near_mem__icache__CAN_FIRE_RL_rl_start_cache_refill &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__EN_req ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_cache_refill_rsps_loop = RTL__near_mem__icache__master_xactor_f_rd_data$EMPTY_N && RTL__near_mem__icache__rg_state ==4'd9; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop = RTL__near_mem__icache__CAN_FIRE_RL_rl_cache_refill_rsps_loop &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__EN_req ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_rereq = RTL__near_mem__icache__rg_state ==4'd10; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq = RTL__near_mem__icache__CAN_FIRE_RL_rl_rereq &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__EN_req ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_ST_AMO_response = RTL__near_mem__icache__rg_state ==4'd11; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_ST_AMO_response = RTL__near_mem__icache__CAN_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_io_read_req = RTL__near_mem__icache__master_xactor_f_rd_addr$FULL_N && RTL__near_mem__icache__rg_state ==4'd12&&! RTL__near_mem__icache__rg_op && RTL__near_mem__icache__b__h14485 ==4'd0; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req = RTL__near_mem__icache__CAN_FIRE_RL_rl_io_read_req &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_io_read_rsp = RTL__near_mem__icache__master_xactor_f_rd_data$EMPTY_N && RTL__near_mem__icache__rg_state ==4'd13; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp = RTL__near_mem__icache__CAN_FIRE_RL_rl_io_read_rsp &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_maintain_io_read_rsp = RTL__near_mem__icache__rg_state ==4'd14; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_maintain_io_read_rsp = RTL__near_mem__icache__CAN_FIRE_RL_rl_maintain_io_read_rsp ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_io_write_req = RTL__near_mem__icache__f_fabric_write_reqs$FULL_N && RTL__near_mem__icache__rg_state ==4'd12&& RTL__near_mem__icache__rg_op ; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req = RTL__near_mem__icache__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_discard_write_rsp = RTL__near_mem__icache__b__h14485 !=4'd0&& RTL__near_mem__icache__master_xactor_f_wr_resp$EMPTY_N ; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp = RTL__near_mem__icache__CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_drive_exception_rsp = RTL__near_mem__icache__rg_state ==4'd4; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_drive_exception_rsp = RTL__near_mem__icache__rg_state ==4'd4; 
  assign  RTL__near_mem__icache__CAN_FIRE_RL_rl_start_reset = RTL__near_mem__icache__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset = RTL__near_mem__icache__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_1 = RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_2 = RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 ; 
  assign  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__SEL_3 = RTL__near_mem__icache__WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL__near_mem__icache__WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__SEL_1 = RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op ; 
  assign  RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 = RTL__near_mem__icache__EN_req && RTL__near_mem__icache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 ; 
  assign  RTL__near_mem__icache__MUX_ram_word64_set$a_put_1__SEL_1 = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2 = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]!=2'd3; 
  assign  RTL__near_mem__icache__MUX_rg_error_during_refill$write_1__SEL_1 = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_1 = RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_2 = RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__SEL_2 = RTL__near_mem__icache__f_reset_reqs$EMPTY_N && RTL__near_mem__icache__rg_state !=4'd1; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__SEL_3 = RTL__near_mem__icache__CAN_FIRE_RL_rl_io_write_req &&! RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__SEL_7 = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]==2'd3; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__SEL_9 = RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 ; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__SEL_10 = RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127; 
  always @(          RTL__near_mem__icache__rg_f3                          or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247                 or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276                or   RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32               or   RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__word64__h5094             or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264            or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285           or   RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  )
         begin 
             case ( RTL__near_mem__icache__rg_f3 )
              3 'b0: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 ;
              3 'b001: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 ;
              3 'b010: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 ;
              3 'b011: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  =( RTL__near_mem__icache__rg_addr [2:0]==3'h0) ?  RTL__near_mem__icache__word64__h5094 :64'd0;
              3 'b100: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 ;
              3 'b101: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 ;
              3 'b110: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  = RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 ;
              3 'd7: 
                  RTL__near_mem__icache__MUX_dw_output_ld_val$wset_1__VAL_2  =64'd0;endcase
         end
  assign  RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__VAL_1 ={ RTL__near_mem__icache__rg_f3 , RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_st_amo_val }; 
  assign  RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__VAL_2 ={ RTL__near_mem__icache__rg_f3 , RTL__near_mem__icache__rg_pa , RTL__near_mem__icache__rg_st_amo_val }; 
  assign  RTL__near_mem__icache__MUX_master_xactor_f_rd_addr$enq_1__VAL_1 ={4'd0, RTL__near_mem__icache__cline_fabric_addr__h14584 ,29'd7143424}; 
  assign  RTL__near_mem__icache__MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ={4'd0, RTL__near_mem__icache__fabric_addr__h17243 ,8'd0, RTL__near_mem__icache__value__h17372 ,18'd65536}; 
  assign  RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ={3'd4, RTL__near_mem__icache__rg_pa [31:12]}; 
  assign  RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_2 = RTL__near_mem__icache__rg_word64_set_in_cache +9'd1; 
  assign  RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_4 ={ RTL__near_mem__icache__rg_addr [11:5],2'd0}; 
  assign  RTL__near_mem__icache__MUX_rg_cset_in_cache$write_1__VAL_1 = RTL__near_mem__icache__rg_cset_in_cache +7'd1; 
  assign  RTL__near_mem__icache__MUX_rg_exc_code$write_1__VAL_1 = RTL__near_mem__icache__req_op  ? 4'd6:4'd4; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__VAL_1 = RTL__near_mem__icache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539  ? 4'd4:4'd3; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__VAL_4 =( RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0) ? 4'd14:4'd4; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__VAL_7 =( RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__icache__rg_error_during_refill ) ? 4'd4:4'd10; 
  assign  RTL__near_mem__icache__MUX_rg_state$write_1__VAL_9 =( RTL__near_mem__icache__dmem_not_imem &&! RTL__near_mem__icache__soc_map$m_is_mem_addr ) ? 4'd12:( RTL__near_mem__icache__rg_op  ? 4'd11:4'd8); 
  assign  RTL__near_mem__icache__dw_valid$whas = RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 || RTL__near_mem__icache__WILL_FIRE_RL_rl_drive_exception_rsp || RTL__near_mem__icache__WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL__near_mem__icache__WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port0__write_1 = RTL__near_mem__icache__ctr_wr_rsps_pending_crg +4'd1; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port1__write_1 = RTL__near_mem__icache__b__h14485 -4'd1; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port2__read = RTL__near_mem__icache__CAN_FIRE_RL_rl_discard_write_rsp  ?  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port1__write_1 : RTL__near_mem__icache__b__h14485 ; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$EN_port2__write = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port3__read = RTL__near_mem__icache__ctr_wr_rsps_pending_crg$EN_port2__write  ? 4'd0: RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port2__read ; 
  assign  RTL__near_mem__icache__cfg_verbosity$D_IN = RTL__near_mem__icache__set_verbosity_verbosity ; 
  assign  RTL__near_mem__icache__cfg_verbosity$EN = RTL__near_mem__icache__EN_set_verbosity ; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$D_IN = RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port3__read ; 
  assign  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$EN =1'b1; 
  assign  RTL__near_mem__icache__rg_addr$D_IN = RTL__near_mem__icache__req_addr ; 
  assign  RTL__near_mem__icache__rg_addr$EN = RTL__near_mem__icache__EN_req ; (* RTL__near_mem__icache__keep *)
    wire[6:0] RTL__near_mem__icache__MUX_rg_cset_in_cache$write_1__VAL_1_any_val ; 
  assign  RTL__near_mem__icache__rg_cset_in_cache$D_IN = RTL__near_mem__icache__WILL_FIRE_RL_rl_reset  ?  RTL__near_mem__icache__MUX_rg_cset_in_cache$write_1__VAL_1_any_val :7'd0; 
  assign  RTL__near_mem__icache__rg_cset_in_cache$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_reset || RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__icache__rg_error_during_refill$D_IN = RTL__near_mem__icache__MUX_rg_error_during_refill$write_1__SEL_1 ; 
  assign  RTL__near_mem__icache__rg_error_during_refill$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill ; 
  always @(      RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_1                  or   RTL__near_mem__icache__MUX_rg_exc_code$write_1__VAL_1             or   RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_2            or   RTL__near_mem__icache__MUX_rg_error_during_refill$write_1__SEL_1           or   RTL__near_mem__icache__access_exc_code__h2256  )
         case (1'b1) 
          RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_1  : 
              RTL__near_mem__icache__rg_exc_code$D_IN  = RTL__near_mem__icache__MUX_rg_exc_code$write_1__VAL_1 ; 
          RTL__near_mem__icache__MUX_rg_exc_code$write_1__SEL_2  : 
              RTL__near_mem__icache__rg_exc_code$D_IN  =4'd5; 
          RTL__near_mem__icache__MUX_rg_error_during_refill$write_1__SEL_1  : 
              RTL__near_mem__icache__rg_exc_code$D_IN  = RTL__near_mem__icache__access_exc_code__h2256 ;
          default : 
              RTL__near_mem__icache__rg_exc_code$D_IN  =4'b1010;endcase
  assign  RTL__near_mem__icache__rg_exc_code$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL__near_mem__icache__rg_f3$D_IN = RTL__near_mem__icache__req_f3 ; 
  assign  RTL__near_mem__icache__rg_f3$EN = RTL__near_mem__icache__EN_req ; 
  assign  RTL__near_mem__icache__rg_ld_val$D_IN = RTL__near_mem__icache__ld_val__h17594 ; 
  assign  RTL__near_mem__icache__rg_ld_val$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp ; 
  assign  RTL__near_mem__icache__rg_lower_word32$D_IN =32'h0; 
  assign  RTL__near_mem__icache__rg_lower_word32$EN =1'b0; 
  assign  RTL__near_mem__icache__rg_lower_word32_full$D_IN =1'd0; 
  assign  RTL__near_mem__icache__rg_lower_word32_full$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL__near_mem__icache__rg_op$D_IN = RTL__near_mem__icache__req_op ; 
  assign  RTL__near_mem__icache__rg_op$EN = RTL__near_mem__icache__EN_req ; 
  assign  RTL__near_mem__icache__rg_pa$D_IN = RTL__near_mem__icache__EN_req  ?  RTL__near_mem__icache__req_addr : RTL__near_mem__icache__rg_addr ; 
  assign  RTL__near_mem__icache__rg_pa$EN = RTL__near_mem__icache__EN_req || RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp ; 
  assign  RTL__near_mem__icache__rg_pte_pa$D_IN =32'h0; 
  assign  RTL__near_mem__icache__rg_pte_pa$EN =1'b0; 
  assign  RTL__near_mem__icache__rg_st_amo_val$D_IN = RTL__near_mem__icache__req_st_value ; 
  assign  RTL__near_mem__icache__rg_st_amo_val$EN = RTL__near_mem__icache__EN_req ; 
  always @(               RTL__near_mem__icache__EN_req                                    or   RTL__near_mem__icache__MUX_rg_state$write_1__VAL_1                      or   RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset                     or   RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req                    or   RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp                   or   RTL__near_mem__icache__MUX_rg_state$write_1__VAL_4                  or   RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req                 or   RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq                or   RTL__near_mem__icache__MUX_rg_state$write_1__SEL_7               or   RTL__near_mem__icache__MUX_rg_state$write_1__VAL_7              or   RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill             or   RTL__near_mem__icache__MUX_rg_state$write_1__SEL_9            or   RTL__near_mem__icache__MUX_rg_state$write_1__VAL_9           or   RTL__near_mem__icache__MUX_rg_state$write_1__SEL_10  )
         case (1'b1) 
          RTL__near_mem__icache__EN_req  : 
              RTL__near_mem__icache__rg_state$D_IN  = RTL__near_mem__icache__MUX_rg_state$write_1__VAL_1 ; 
          RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset  : 
              RTL__near_mem__icache__rg_state$D_IN  =4'd1; 
          RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req  : 
              RTL__near_mem__icache__rg_state$D_IN  =4'd11; 
          RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp  : 
              RTL__near_mem__icache__rg_state$D_IN  = RTL__near_mem__icache__MUX_rg_state$write_1__VAL_4 ; 
          RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req  : 
              RTL__near_mem__icache__rg_state$D_IN  =4'd13; 
          RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq  : 
              RTL__near_mem__icache__rg_state$D_IN  =4'd3; 
          RTL__near_mem__icache__MUX_rg_state$write_1__SEL_7  : 
              RTL__near_mem__icache__rg_state$D_IN  = RTL__near_mem__icache__MUX_rg_state$write_1__VAL_7 ; 
          RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  : 
              RTL__near_mem__icache__rg_state$D_IN  =4'd9; 
          RTL__near_mem__icache__MUX_rg_state$write_1__SEL_9  : 
              RTL__near_mem__icache__rg_state$D_IN  = RTL__near_mem__icache__MUX_rg_state$write_1__VAL_9 ; 
          RTL__near_mem__icache__MUX_rg_state$write_1__SEL_10  : 
              RTL__near_mem__icache__rg_state$D_IN  =4'd2;
          default : 
              RTL__near_mem__icache__rg_state$D_IN  =4'b1010;endcase
  assign  RTL__near_mem__icache__rg_state$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127|| RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]==2'd3|| RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 || RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp || RTL__near_mem__icache__EN_req || RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset || RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq || RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req || RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL__near_mem__icache__rg_word64_set_in_cache$D_IN = RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2  ?  RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_2 : RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_4 ; 
  assign  RTL__near_mem__icache__rg_word64_set_in_cache$EN = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]!=2'd3|| RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs$D_IN = RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__SEL_1  ?  RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__VAL_1 : RTL__near_mem__icache__MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs$ENQ = RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op || RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs$DEQ = RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__icache__f_fabric_write_reqs$CLR =1'b0; 
  assign  RTL__near_mem__icache__f_reset_reqs$D_IN =! RTL__near_mem__icache__EN_server_reset_request_put ; 
  assign  RTL__near_mem__icache__f_reset_reqs$ENQ = RTL__near_mem__icache__EN_server_reset_request_put || RTL__near_mem__icache__EN_server_flush_request_put ; 
  assign  RTL__near_mem__icache__f_reset_reqs$DEQ = RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127; 
  assign  RTL__near_mem__icache__f_reset_reqs$CLR =1'b0; 
  assign  RTL__near_mem__icache__f_reset_rsps$D_IN = RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__f_reset_rsps$ENQ = RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127; 
  assign  RTL__near_mem__icache__f_reset_rsps$DEQ = RTL__near_mem__icache__EN_server_flush_response_get || RTL__near_mem__icache__EN_server_reset_response_get ; 
  assign  RTL__near_mem__icache__f_reset_rsps$CLR =1'b0; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr$D_IN = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  ?  RTL__near_mem__icache__MUX_master_xactor_f_rd_addr$enq_1__VAL_1 : RTL__near_mem__icache__MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr$ENQ = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr$DEQ = RTL__near_mem__icache__master_xactor_f_rd_addr$EMPTY_N && RTL__near_mem__icache__mem_master_arready ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_addr$CLR = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data$D_IN ={ RTL__near_mem__icache__mem_master_rid , RTL__near_mem__icache__mem_master_rdata , RTL__near_mem__icache__mem_master_rresp , RTL__near_mem__icache__mem_master_rlast }; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data$ENQ = RTL__near_mem__icache__mem_master_rvalid && RTL__near_mem__icache__master_xactor_f_rd_data$FULL_N ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data$DEQ = RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp || RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop ; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_data$CLR = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr$D_IN ={4'd0, RTL__near_mem__icache__mem_req_wr_addr_awaddr__h2473 ,8'd0, RTL__near_mem__icache__x__h2520 ,18'd65536}; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr$ENQ = RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr$DEQ = RTL__near_mem__icache__master_xactor_f_wr_addr$EMPTY_N && RTL__near_mem__icache__mem_master_awready ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_addr$CLR = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data$D_IN ={ RTL__near_mem__icache__mem_req_wr_data_wdata__h2699 , RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700 ,1'd1}; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data$ENQ = RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data$DEQ = RTL__near_mem__icache__master_xactor_f_wr_data$EMPTY_N && RTL__near_mem__icache__mem_master_wready ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_data$CLR = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp$D_IN ={ RTL__near_mem__icache__mem_master_bid , RTL__near_mem__icache__mem_master_bresp }; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp$ENQ = RTL__near_mem__icache__mem_master_bvalid && RTL__near_mem__icache__master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp$DEQ = RTL__near_mem__icache__CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL__near_mem__icache__master_xactor_f_wr_resp$CLR = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset &&! RTL__near_mem__icache__f_reset_reqs$D_OUT ; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$ADDRA = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  ?  RTL__near_mem__icache__rg_addr [11:5]: RTL__near_mem__icache__rg_cset_in_cache ; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$ADDRB = RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ?  RTL__near_mem__icache__req_addr [11:5]: RTL__near_mem__icache__rg_addr [11:5]; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$DIA = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  ?  RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 :23'd2796202; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$DIB = RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ? 23'b01010101010101010101010:23'b01010101010101010101010; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$WEA =1'd1; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$WEB =1'd0; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$ENA = RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill || RTL__near_mem__icache__WILL_FIRE_RL_rl_reset ; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset$ENB = RTL__near_mem__icache__EN_req && RTL__near_mem__icache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq ; 
  assign  RTL__near_mem__icache__ram_word64_set$ADDRA = RTL__near_mem__icache__MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL__near_mem__icache__rg_word64_set_in_cache : RTL__near_mem__icache__rg_addr [11:3]; 
  always @(         RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                        or   RTL__near_mem__icache__req_addr                or   RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2               or   RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_2              or   RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq             or   RTL__near_mem__icache__rg_addr            or   RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill           or   RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_4  )
         begin 
             case (1'b1) 
              RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL__near_mem__icache__ram_word64_set$ADDRB  = RTL__near_mem__icache__req_addr [11:3]; 
              RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL__near_mem__icache__ram_word64_set$ADDRB  = RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_2 ; 
              RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq  : 
                  RTL__near_mem__icache__ram_word64_set$ADDRB  = RTL__near_mem__icache__rg_addr [11:3]; 
              RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL__near_mem__icache__ram_word64_set$ADDRB  = RTL__near_mem__icache__MUX_ram_word64_set$b_put_2__VAL_4 ;
              default : 
                  RTL__near_mem__icache__ram_word64_set$ADDRB  =9'b010101010;endcase
         end
  assign  RTL__near_mem__icache__ram_word64_set$DIA = RTL__near_mem__icache__MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:3]: RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 ; 
  always @(     RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                or   RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2            or   RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq           or   RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  )
         begin 
             case (1'b1) 
              RTL__near_mem__icache__MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL__near_mem__icache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL__near_mem__icache__MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL__near_mem__icache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq  : 
                  RTL__near_mem__icache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL__near_mem__icache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;
              default : 
                  RTL__near_mem__icache__ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL__near_mem__icache__ram_word64_set$WEA =1'd1; 
  assign  RTL__near_mem__icache__ram_word64_set$WEB =1'd0; 
  assign  RTL__near_mem__icache__ram_word64_set$ENA = RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 ; 
  assign  RTL__near_mem__icache__ram_word64_set$ENB = RTL__near_mem__icache__EN_req && RTL__near_mem__icache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]!=2'd3|| RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq || RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL__near_mem__icache__soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL__near_mem__icache__soc_map$m_is_mem_addr_addr ={32'd0, RTL__near_mem__icache__rg_addr }; 
  assign  RTL__near_mem__icache__soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 = RTL__near_mem__icache__cfg_verbosity >4'd1; 
  assign  RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 = RTL__near_mem__icache__cfg_verbosity >4'd2; 
  assign  RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 =(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op && RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL__near_mem__icache__NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 =(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&&! RTL__near_mem__icache__rg_op && RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL__near_mem__icache__NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 = RTL__near_mem__icache__req_f3 [1:0]!=2'b0&&( RTL__near_mem__icache__req_f3 [1:0]!=2'b01|| RTL__near_mem__icache__req_addr [0])&&( RTL__near_mem__icache__req_f3 [1:0]!=2'b10|| RTL__near_mem__icache__req_addr [1:0]!=2'b0)&&( RTL__near_mem__icache__req_f3 [1:0]!=2'b11|| RTL__near_mem__icache__req_addr [2:0]!=3'b0); 
  assign  RTL__near_mem__icache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 =! RTL__near_mem__icache__rg_op && RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL__near_mem__icache___theResult___snd_fst__h2707 = RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [63:0]<< RTL__near_mem__icache__shift_bits__h2487 ; 
  assign  RTL__near_mem__icache__access_exc_code__h2256 = RTL__near_mem__icache__dmem_not_imem  ? ( RTL__near_mem__icache__rg_op  ? 4'd7:4'd5):4'd1; 
  assign  RTL__near_mem__icache__b__h14485 = RTL__near_mem__icache__CAN_FIRE_RL_rl_fabric_send_write_req  ?  RTL__near_mem__icache__ctr_wr_rsps_pending_crg$port0__write_1 : RTL__near_mem__icache__ctr_wr_rsps_pending_crg ; 
  assign  RTL__near_mem__icache__cline_addr__h14583 ={ RTL__near_mem__icache__rg_pa [31:5],5'd0}; 
  assign  RTL__near_mem__icache__cline_fabric_addr__h14584 ={32'd0, RTL__near_mem__icache__cline_addr__h14583 }; 
  assign  RTL__near_mem__icache__dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 = RTL__near_mem__icache__dmem_not_imem &&! RTL__near_mem__icache__soc_map$m_is_mem_addr || RTL__near_mem__icache__rg_op ||! RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]||! RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL__near_mem__icache__fabric_addr__h17243 ={32'd0, RTL__near_mem__icache__rg_pa }; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [10:3]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [18:11]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [18:3]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [26:19]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [34:19]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [34:27]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [34:3]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [42:35]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [50:35]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [50:43]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [58:51]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:35]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:51]; 
  assign  RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 = RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:59]; 
  assign  RTL__near_mem__icache__mem_req_wr_addr_awaddr__h2473 ={32'd0, RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [95:64]}; 
  assign  RTL__near_mem__icache__pa_ctag__h4952 ={2'd0, RTL__near_mem__icache__rg_addr [31:12]}; 
  assign  RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 = RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [21:0]== RTL__near_mem__icache__pa_ctag__h4952 ; 
  assign  RTL__near_mem__icache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 = RTL__near_mem__icache__req_f3 [1:0]==2'b0|| RTL__near_mem__icache__req_f3 [1:0]==2'b01&&! RTL__near_mem__icache__req_addr [0]|| RTL__near_mem__icache__req_f3 [1:0]==2'b10&& RTL__near_mem__icache__req_addr [1:0]==2'b0|| RTL__near_mem__icache__req_f3 [1:0]==2'b11&& RTL__near_mem__icache__req_addr [2:0]==3'b0; 
  assign  RTL__near_mem__icache__result__h11657 ={{56{ RTL__near_mem__icache__word64094_BITS_15_TO_8__q18 [7]}}, RTL__near_mem__icache__word64094_BITS_15_TO_8__q18 }; 
  assign  RTL__near_mem__icache__result__h11685 ={{56{ RTL__near_mem__icache__word64094_BITS_23_TO_16__q19 [7]}}, RTL__near_mem__icache__word64094_BITS_23_TO_16__q19 }; 
  assign  RTL__near_mem__icache__result__h11713 ={{56{ RTL__near_mem__icache__word64094_BITS_31_TO_24__q21 [7]}}, RTL__near_mem__icache__word64094_BITS_31_TO_24__q21 }; 
  assign  RTL__near_mem__icache__result__h11741 ={{56{ RTL__near_mem__icache__word64094_BITS_39_TO_32__q22 [7]}}, RTL__near_mem__icache__word64094_BITS_39_TO_32__q22 }; 
  assign  RTL__near_mem__icache__result__h11769 ={{56{ RTL__near_mem__icache__word64094_BITS_47_TO_40__q25 [7]}}, RTL__near_mem__icache__word64094_BITS_47_TO_40__q25 }; 
  assign  RTL__near_mem__icache__result__h11797 ={{56{ RTL__near_mem__icache__word64094_BITS_55_TO_48__q26 [7]}}, RTL__near_mem__icache__word64094_BITS_55_TO_48__q26 }; 
  assign  RTL__near_mem__icache__result__h11825 ={{56{ RTL__near_mem__icache__word64094_BITS_63_TO_56__q28 [7]}}, RTL__near_mem__icache__word64094_BITS_63_TO_56__q28 }; 
  assign  RTL__near_mem__icache__result__h11870 ={56'd0, RTL__near_mem__icache__word64__h5094 [7:0]}; 
  assign  RTL__near_mem__icache__result__h11898 ={56'd0, RTL__near_mem__icache__word64__h5094 [15:8]}; 
  assign  RTL__near_mem__icache__result__h11926 ={56'd0, RTL__near_mem__icache__word64__h5094 [23:16]}; 
  assign  RTL__near_mem__icache__result__h11954 ={56'd0, RTL__near_mem__icache__word64__h5094 [31:24]}; 
  assign  RTL__near_mem__icache__result__h11982 ={56'd0, RTL__near_mem__icache__word64__h5094 [39:32]}; 
  assign  RTL__near_mem__icache__result__h12010 ={56'd0, RTL__near_mem__icache__word64__h5094 [47:40]}; 
  assign  RTL__near_mem__icache__result__h12038 ={56'd0, RTL__near_mem__icache__word64__h5094 [55:48]}; 
  assign  RTL__near_mem__icache__result__h12066 ={56'd0, RTL__near_mem__icache__word64__h5094 [63:56]}; 
  assign  RTL__near_mem__icache__result__h12111 ={{48{ RTL__near_mem__icache__word64094_BITS_15_TO_0__q16 [15]}}, RTL__near_mem__icache__word64094_BITS_15_TO_0__q16 }; 
  assign  RTL__near_mem__icache__result__h12139 ={{48{ RTL__near_mem__icache__word64094_BITS_31_TO_16__q20 [15]}}, RTL__near_mem__icache__word64094_BITS_31_TO_16__q20 }; 
  assign  RTL__near_mem__icache__result__h12167 ={{48{ RTL__near_mem__icache__word64094_BITS_47_TO_32__q23 [15]}}, RTL__near_mem__icache__word64094_BITS_47_TO_32__q23 }; 
  assign  RTL__near_mem__icache__result__h12195 ={{48{ RTL__near_mem__icache__word64094_BITS_63_TO_48__q27 [15]}}, RTL__near_mem__icache__word64094_BITS_63_TO_48__q27 }; 
  assign  RTL__near_mem__icache__result__h12236 ={48'd0, RTL__near_mem__icache__word64__h5094 [15:0]}; 
  assign  RTL__near_mem__icache__result__h12264 ={48'd0, RTL__near_mem__icache__word64__h5094 [31:16]}; 
  assign  RTL__near_mem__icache__result__h12292 ={48'd0, RTL__near_mem__icache__word64__h5094 [47:32]}; 
  assign  RTL__near_mem__icache__result__h12320 ={48'd0, RTL__near_mem__icache__word64__h5094 [63:48]}; 
  assign  RTL__near_mem__icache__result__h12361 ={{32{ RTL__near_mem__icache__word64094_BITS_31_TO_0__q17 [31]}}, RTL__near_mem__icache__word64094_BITS_31_TO_0__q17 }; 
  assign  RTL__near_mem__icache__result__h12389 ={{32{ RTL__near_mem__icache__word64094_BITS_63_TO_32__q24 [31]}}, RTL__near_mem__icache__word64094_BITS_63_TO_32__q24 }; 
  assign  RTL__near_mem__icache__result__h12428 ={32'd0, RTL__near_mem__icache__word64__h5094 [31:0]}; 
  assign  RTL__near_mem__icache__result__h12456 ={32'd0, RTL__near_mem__icache__word64__h5094 [63:32]}; 
  assign  RTL__near_mem__icache__result__h17654 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 }; 
  assign  RTL__near_mem__icache__result__h17684 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 }; 
  assign  RTL__near_mem__icache__result__h17711 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 }; 
  assign  RTL__near_mem__icache__result__h17738 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 }; 
  assign  RTL__near_mem__icache__result__h17765 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 }; 
  assign  RTL__near_mem__icache__result__h17792 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 }; 
  assign  RTL__near_mem__icache__result__h17819 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 }; 
  assign  RTL__near_mem__icache__result__h17846 ={{56{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 [7]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 }; 
  assign  RTL__near_mem__icache__result__h17890 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [10:3]}; 
  assign  RTL__near_mem__icache__result__h17917 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [18:11]}; 
  assign  RTL__near_mem__icache__result__h17944 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [26:19]}; 
  assign  RTL__near_mem__icache__result__h17971 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [34:27]}; 
  assign  RTL__near_mem__icache__result__h17998 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [42:35]}; 
  assign  RTL__near_mem__icache__result__h18025 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [50:43]}; 
  assign  RTL__near_mem__icache__result__h18052 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [58:51]}; 
  assign  RTL__near_mem__icache__result__h18079 ={56'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:59]}; 
  assign  RTL__near_mem__icache__result__h18123 ={{48{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 [15]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 }; 
  assign  RTL__near_mem__icache__result__h18150 ={{48{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 [15]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 }; 
  assign  RTL__near_mem__icache__result__h18177 ={{48{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 [15]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 }; 
  assign  RTL__near_mem__icache__result__h18204 ={{48{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 [15]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 }; 
  assign  RTL__near_mem__icache__result__h18244 ={48'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [18:3]}; 
  assign  RTL__near_mem__icache__result__h18271 ={48'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [34:19]}; 
  assign  RTL__near_mem__icache__result__h18298 ={48'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [50:35]}; 
  assign  RTL__near_mem__icache__result__h18325 ={48'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:51]}; 
  assign  RTL__near_mem__icache__result__h18365 ={{32{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 [31]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 }; 
  assign  RTL__near_mem__icache__result__h18392 ={{32{ RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 [31]}}, RTL__near_mem__icache__master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 }; 
  assign  RTL__near_mem__icache__result__h18430 ={32'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [34:3]}; 
  assign  RTL__near_mem__icache__result__h18457 ={32'd0, RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:35]}; 
  assign  RTL__near_mem__icache__result__h5301 ={{56{ RTL__near_mem__icache__word64094_BITS_7_TO_0__q15 [7]}}, RTL__near_mem__icache__word64094_BITS_7_TO_0__q15 }; 
  assign  RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 = RTL__near_mem__icache__rg_op && RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL__near_mem__icache__shift_bits__h2487 ={ RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [66:64],3'b0}; 
  assign  RTL__near_mem__icache__strobe64__h2637 =8'b00000001<< RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL__near_mem__icache__strobe64__h2639 =8'b00000011<< RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL__near_mem__icache__strobe64__h2641 =8'b00001111<< RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL__near_mem__icache__word64094_BITS_15_TO_0__q16 = RTL__near_mem__icache__word64__h5094 [15:0]; 
  assign  RTL__near_mem__icache__word64094_BITS_15_TO_8__q18 = RTL__near_mem__icache__word64__h5094 [15:8]; 
  assign  RTL__near_mem__icache__word64094_BITS_23_TO_16__q19 = RTL__near_mem__icache__word64__h5094 [23:16]; 
  assign  RTL__near_mem__icache__word64094_BITS_31_TO_0__q17 = RTL__near_mem__icache__word64__h5094 [31:0]; 
  assign  RTL__near_mem__icache__word64094_BITS_31_TO_16__q20 = RTL__near_mem__icache__word64__h5094 [31:16]; 
  assign  RTL__near_mem__icache__word64094_BITS_31_TO_24__q21 = RTL__near_mem__icache__word64__h5094 [31:24]; 
  assign  RTL__near_mem__icache__word64094_BITS_39_TO_32__q22 = RTL__near_mem__icache__word64__h5094 [39:32]; 
  assign  RTL__near_mem__icache__word64094_BITS_47_TO_32__q23 = RTL__near_mem__icache__word64__h5094 [47:32]; 
  assign  RTL__near_mem__icache__word64094_BITS_47_TO_40__q25 = RTL__near_mem__icache__word64__h5094 [47:40]; 
  assign  RTL__near_mem__icache__word64094_BITS_55_TO_48__q26 = RTL__near_mem__icache__word64__h5094 [55:48]; 
  assign  RTL__near_mem__icache__word64094_BITS_63_TO_32__q24 = RTL__near_mem__icache__word64__h5094 [63:32]; 
  assign  RTL__near_mem__icache__word64094_BITS_63_TO_48__q27 = RTL__near_mem__icache__word64__h5094 [63:48]; 
  assign  RTL__near_mem__icache__word64094_BITS_63_TO_56__q28 = RTL__near_mem__icache__word64__h5094 [63:56]; 
  assign  RTL__near_mem__icache__word64094_BITS_7_TO_0__q15 = RTL__near_mem__icache__word64__h5094 [7:0]; 
  assign  RTL__near_mem__icache__word64__h5094 = RTL__near_mem__icache__ram_word64_set$DOB & RTL__near_mem__icache__y__h5337 ; 
  assign  RTL__near_mem__icache__y__h5337 ={64{ RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]&& RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 }}; 
  always @(  RTL__near_mem__icache__f_fabric_write_reqs$D_OUT  )
         begin 
             case ( RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL__near_mem__icache__x__h2520  =3'b0;
              2 'b01: 
                  RTL__near_mem__icache__x__h2520  =3'b001;
              2 'b10: 
                  RTL__near_mem__icache__x__h2520  =3'b010;
              2 'b11: 
                  RTL__near_mem__icache__x__h2520  =3'b011;endcase
         end
  always @(  RTL__near_mem__icache__rg_f3  )
         begin 
             case ( RTL__near_mem__icache__rg_f3 [1:0])
              2 'b0: 
                  RTL__near_mem__icache__value__h17372  =3'b0;
              2 'b01: 
                  RTL__near_mem__icache__value__h17372  =3'b001;
              2 'b10: 
                  RTL__near_mem__icache__value__h17372  =3'b010;
              2 'd3: 
                  RTL__near_mem__icache__value__h17372  =3'b011;endcase
         end
  always @(     RTL__near_mem__icache__f_fabric_write_reqs$D_OUT                or   RTL__near_mem__icache__strobe64__h2637            or   RTL__near_mem__icache__strobe64__h2639           or   RTL__near_mem__icache__strobe64__h2641  )
         begin 
             case ( RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700  = RTL__near_mem__icache__strobe64__h2637 ;
              2 'b01: 
                  RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700  = RTL__near_mem__icache__strobe64__h2639 ;
              2 'b10: 
                  RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700  = RTL__near_mem__icache__strobe64__h2641 ;
              2 'b11: 
                  RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700  =8'b11111111;endcase
         end
  always @(   RTL__near_mem__icache__f_fabric_write_reqs$D_OUT            or   RTL__near_mem__icache___theResult___snd_fst__h2707  )
         begin 
             case ( RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [97:96])
              2 'b0,2'b01,2'b10: 
                  RTL__near_mem__icache__mem_req_wr_data_wdata__h2699  = RTL__near_mem__icache___theResult___snd_fst__h2707 ;
              2 'd3: 
                  RTL__near_mem__icache__mem_req_wr_data_wdata__h2699  = RTL__near_mem__icache__f_fabric_write_reqs$D_OUT [63:0];endcase
         end
  always @(      RTL__near_mem__icache__rg_addr                  or   RTL__near_mem__icache__result__h12111             or   RTL__near_mem__icache__result__h12139            or   RTL__near_mem__icache__result__h12167           or   RTL__near_mem__icache__result__h12195  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__icache__result__h12111 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__icache__result__h12139 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__icache__result__h12167 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL__near_mem__icache__result__h12195 ;
              default : 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  =64'd0;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__ram_word64_set$DOB           or   RTL__near_mem__icache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:16], RTL__near_mem__icache__rg_st_amo_val [15:0]};
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:32], RTL__near_mem__icache__rg_st_amo_val [15:0], RTL__near_mem__icache__ram_word64_set$DOB [15:0]};
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:48], RTL__near_mem__icache__rg_st_amo_val [15:0], RTL__near_mem__icache__ram_word64_set$DOB [31:0]};
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL__near_mem__icache__rg_st_amo_val [15:0], RTL__near_mem__icache__ram_word64_set$DOB [47:0]};
              default : 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  = RTL__near_mem__icache__ram_word64_set$DOB ;endcase
         end
  always @(          RTL__near_mem__icache__rg_addr                          or   RTL__near_mem__icache__result__h5301                 or   RTL__near_mem__icache__result__h11657                or   RTL__near_mem__icache__result__h11685               or   RTL__near_mem__icache__result__h11713              or   RTL__near_mem__icache__result__h11741             or   RTL__near_mem__icache__result__h11769            or   RTL__near_mem__icache__result__h11797           or   RTL__near_mem__icache__result__h11825  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h5301 ;
              3 'h1: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11657 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11685 ;
              3 'h3: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11713 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11741 ;
              3 'h5: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11769 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11797 ;
              3 'h7: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL__near_mem__icache__result__h11825 ;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__ram_word64_set$DOB           or   RTL__near_mem__icache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:8], RTL__near_mem__icache__rg_st_amo_val [7:0]};
              3 'h1: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:16], RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [7:0]};
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:24], RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [15:0]};
              3 'h3: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:32], RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [23:0]};
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:40], RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [31:0]};
              3 'h5: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:48], RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [39:0]};
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:56], RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [47:0]};
              3 'h7: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL__near_mem__icache__rg_st_amo_val [7:0], RTL__near_mem__icache__ram_word64_set$DOB [55:0]};endcase
         end
  always @(      RTL__near_mem__icache__rg_addr                  or   RTL__near_mem__icache__result__h18244             or   RTL__near_mem__icache__result__h18271            or   RTL__near_mem__icache__result__h18298           or   RTL__near_mem__icache__result__h18325  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__icache__result__h18244 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__icache__result__h18271 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__icache__result__h18298 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL__near_mem__icache__result__h18325 ;
              default : 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  =64'd0;endcase
         end
  always @(      RTL__near_mem__icache__rg_addr                  or   RTL__near_mem__icache__result__h12236             or   RTL__near_mem__icache__result__h12264            or   RTL__near_mem__icache__result__h12292           or   RTL__near_mem__icache__result__h12320  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__icache__result__h12236 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__icache__result__h12264 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__icache__result__h12292 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL__near_mem__icache__result__h12320 ;
              default : 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  =64'd0;endcase
         end
  always @(      RTL__near_mem__icache__rg_addr                  or   RTL__near_mem__icache__result__h18123             or   RTL__near_mem__icache__result__h18150            or   RTL__near_mem__icache__result__h18177           or   RTL__near_mem__icache__result__h18204  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__icache__result__h18123 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__icache__result__h18150 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__icache__result__h18177 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL__near_mem__icache__result__h18204 ;
              default : 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  =64'd0;endcase
         end
  always @(          RTL__near_mem__icache__rg_addr                          or   RTL__near_mem__icache__result__h17890                 or   RTL__near_mem__icache__result__h17917                or   RTL__near_mem__icache__result__h17944               or   RTL__near_mem__icache__result__h17971              or   RTL__near_mem__icache__result__h17998             or   RTL__near_mem__icache__result__h18025            or   RTL__near_mem__icache__result__h18052           or   RTL__near_mem__icache__result__h18079  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h17890 ;
              3 'h1: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h17917 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h17944 ;
              3 'h3: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h17971 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h17998 ;
              3 'h5: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h18025 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h18052 ;
              3 'h7: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL__near_mem__icache__result__h18079 ;endcase
         end
  always @(          RTL__near_mem__icache__rg_addr                          or   RTL__near_mem__icache__result__h11870                 or   RTL__near_mem__icache__result__h11898                or   RTL__near_mem__icache__result__h11926               or   RTL__near_mem__icache__result__h11954              or   RTL__near_mem__icache__result__h11982             or   RTL__near_mem__icache__result__h12010            or   RTL__near_mem__icache__result__h12038           or   RTL__near_mem__icache__result__h12066  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h11870 ;
              3 'h1: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h11898 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h11926 ;
              3 'h3: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h11954 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h11982 ;
              3 'h5: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h12010 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h12038 ;
              3 'h7: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL__near_mem__icache__result__h12066 ;endcase
         end
  always @(          RTL__near_mem__icache__rg_addr                          or   RTL__near_mem__icache__result__h17654                 or   RTL__near_mem__icache__result__h17684                or   RTL__near_mem__icache__result__h17711               or   RTL__near_mem__icache__result__h17738              or   RTL__near_mem__icache__result__h17765             or   RTL__near_mem__icache__result__h17792            or   RTL__near_mem__icache__result__h17819           or   RTL__near_mem__icache__result__h17846  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17654 ;
              3 'h1: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17684 ;
              3 'h2: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17711 ;
              3 'h3: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17738 ;
              3 'h4: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17765 ;
              3 'h5: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17792 ;
              3 'h6: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17819 ;
              3 'h7: 
                  RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL__near_mem__icache__result__h17846 ;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__result__h18365           or   RTL__near_mem__icache__result__h18392  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL__near_mem__icache__result__h18365 ;
              3 'h4: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL__near_mem__icache__result__h18392 ;
              default : 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  =64'd0;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__result__h18430           or   RTL__near_mem__icache__result__h18457  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL__near_mem__icache__result__h18430 ;
              3 'h4: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL__near_mem__icache__result__h18457 ;
              default : 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  =64'd0;endcase
         end
  always @(          RTL__near_mem__icache__rg_f3                          or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411                 or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439                or   RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29               or   RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT             or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427            or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447           or   RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  )
         begin 
             case ( RTL__near_mem__icache__rg_f3 )
              3 'b0: 
                  RTL__near_mem__icache__ld_val__h17594  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 ;
              3 'b001: 
                  RTL__near_mem__icache__ld_val__h17594  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 ;
              3 'b010: 
                  RTL__near_mem__icache__ld_val__h17594  = RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 ;
              3 'b011: 
                  RTL__near_mem__icache__ld_val__h17594  =( RTL__near_mem__icache__rg_addr [2:0]==3'h0) ?  RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:3]:64'd0;
              3 'b100: 
                  RTL__near_mem__icache__ld_val__h17594  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 ;
              3 'b101: 
                  RTL__near_mem__icache__ld_val__h17594  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 ;
              3 'b110: 
                  RTL__near_mem__icache__ld_val__h17594  = RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 ;
              3 'd7: 
                  RTL__near_mem__icache__ld_val__h17594  =64'd0;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__ram_word64_set$DOB           or   RTL__near_mem__icache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL__near_mem__icache__ram_word64_set$DOB [63:32], RTL__near_mem__icache__rg_st_amo_val [31:0]};
              3 'h4: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL__near_mem__icache__rg_st_amo_val [31:0], RTL__near_mem__icache__ram_word64_set$DOB [31:0]};
              default : 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  = RTL__near_mem__icache__ram_word64_set$DOB ;endcase
         end
  always @(       RTL__near_mem__icache__rg_f3                    or   RTL__near_mem__icache__ram_word64_set$DOB              or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157             or   RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167            or   RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31           or   RTL__near_mem__icache__rg_st_amo_val  )
         begin 
             case ( RTL__near_mem__icache__rg_f3 )
              3 'b0: 
                  RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 ;
              3 'b001: 
                  RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__icache__IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 ;
              3 'b010: 
                  RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 ;
              3 'b011: 
                  RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__icache__rg_st_amo_val ;
              default : 
                  RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL__near_mem__icache__ram_word64_set$DOB ;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__result__h12361           or   RTL__near_mem__icache__result__h12389  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL__near_mem__icache__result__h12361 ;
              3 'h4: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL__near_mem__icache__result__h12389 ;
              default : 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  =64'd0;endcase
         end
  always @(    RTL__near_mem__icache__rg_addr              or   RTL__near_mem__icache__result__h12428           or   RTL__near_mem__icache__result__h12456  )
         begin 
             case ( RTL__near_mem__icache__rg_addr [2:0])
              3 'h0: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL__near_mem__icache__result__h12428 ;
              3 'h4: 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL__near_mem__icache__result__h12456 ;
              default : 
                  RTL__near_mem__icache__CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  =64'd0;endcase
         end
  always @( posedge  RTL__near_mem__icache__CLK )
         begin 
             if ( RTL__near_mem__icache__RST_N ==1'b0)
                 begin  
                     RTL__near_mem__icache__cfg_verbosity  <=4'd0; 
                     RTL__near_mem__icache__ctr_wr_rsps_pending_crg  <=4'd0; 
                     RTL__near_mem__icache__rg_cset_in_cache  <=7'd0; 
                     RTL__near_mem__icache__rg_lower_word32_full  <=1'd0; 
                     RTL__near_mem__icache__rg_state  <=4'd0;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__icache__cfg_verbosity$EN ) 
                         RTL__near_mem__icache__cfg_verbosity  <= RTL__near_mem__icache__cfg_verbosity$D_IN ;
                     if ( RTL__near_mem__icache__ctr_wr_rsps_pending_crg$EN ) 
                         RTL__near_mem__icache__ctr_wr_rsps_pending_crg  <= RTL__near_mem__icache__ctr_wr_rsps_pending_crg$D_IN ;
                     if ( RTL__near_mem__icache__rg_cset_in_cache$EN ) 
                         RTL__near_mem__icache__rg_cset_in_cache  <= RTL__near_mem__icache__rg_cset_in_cache$D_IN ;
                     if ( RTL__near_mem__icache__rg_lower_word32_full$EN ) 
                         RTL__near_mem__icache__rg_lower_word32_full  <= RTL__near_mem__icache__rg_lower_word32_full$D_IN ;
                     if ( RTL__near_mem__icache__rg_state$EN ) 
                         RTL__near_mem__icache__rg_state  <= RTL__near_mem__icache__rg_state$D_IN ;
                 end 
             if ( RTL__near_mem__icache__rg_addr$EN ) 
                 RTL__near_mem__icache__rg_addr  <= RTL__near_mem__icache__rg_addr$D_IN ;
             if ( RTL__near_mem__icache__rg_error_during_refill$EN ) 
                 RTL__near_mem__icache__rg_error_during_refill  <= RTL__near_mem__icache__rg_error_during_refill$D_IN ;
             if ( RTL__near_mem__icache__rg_exc_code$EN ) 
                 RTL__near_mem__icache__rg_exc_code  <= RTL__near_mem__icache__rg_exc_code$D_IN ;
             if ( RTL__near_mem__icache__rg_f3$EN ) 
                 RTL__near_mem__icache__rg_f3  <= RTL__near_mem__icache__rg_f3$D_IN ;
             if ( RTL__near_mem__icache__rg_ld_val$EN ) 
                 RTL__near_mem__icache__rg_ld_val  <= RTL__near_mem__icache__rg_ld_val$D_IN ;
             if ( RTL__near_mem__icache__rg_lower_word32$EN ) 
                 RTL__near_mem__icache__rg_lower_word32  <= RTL__near_mem__icache__rg_lower_word32$D_IN ;
             if ( RTL__near_mem__icache__rg_op$EN ) 
                 RTL__near_mem__icache__rg_op  <= RTL__near_mem__icache__rg_op$D_IN ;
             if ( RTL__near_mem__icache__rg_pa$EN ) 
                 RTL__near_mem__icache__rg_pa  <= RTL__near_mem__icache__rg_pa$D_IN ;
             if ( RTL__near_mem__icache__rg_pte_pa$EN ) 
                 RTL__near_mem__icache__rg_pte_pa  <= RTL__near_mem__icache__rg_pte_pa$D_IN ;
             if ( RTL__near_mem__icache__rg_st_amo_val$EN ) 
                 RTL__near_mem__icache__rg_st_amo_val  <= RTL__near_mem__icache__rg_st_amo_val$D_IN ;
             if ( RTL__near_mem__icache__rg_word64_set_in_cache$EN ) 
                 RTL__near_mem__icache__rg_word64_set_in_cache  <= RTL__near_mem__icache__rg_word64_set_in_cache$D_IN ;
         end
  always @( negedge  RTL__near_mem__icache__CLK )
         begin #0;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__ctr_wr_rsps_pending_crg ==4'd15)
                     begin  
                         RTL__near_mem__icache__v__h2948  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h2942  = RTL__near_mem__icache__v__h2948 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__ctr_wr_rsps_pending_crg ==4'd15)$display("%0d: ERROR: CreditCounter: overflow", RTL__near_mem__icache__v__h2942 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__ctr_wr_rsps_pending_crg ==4'd15)$finish(32'd1);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Addr { ","awid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awaddr: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__mem_req_wr_addr_awaddr__h2473 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlen: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awsize: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__x__h2520 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awburst: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlock: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awcache: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awprot: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awqos: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awregion: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awuser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("                       ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Data { ","wdata: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__mem_req_wr_data_wdata__h2699 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wstrb: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__mem_req_wr_data_wstrb__h2700 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wlast: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("True");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wuser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_fabric_send_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127&& RTL__near_mem__icache__cfg_verbosity !=4'd0&&! RTL__near_mem__icache__f_reset_reqs$D_OUT )
                     begin  
                         RTL__near_mem__icache__v__h3848  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h3842  = RTL__near_mem__icache__v__h3848 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127&& RTL__near_mem__icache__cfg_verbosity !=4'd0&&! RTL__near_mem__icache__f_reset_reqs$D_OUT )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL__near_mem__icache__v__h3842 ,"D_MMU_Cache",$signed(32'd128),$signed(32'd1));
                      else $display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL__near_mem__icache__v__h3842 ,"I_MMU_Cache",$signed(32'd128),$signed(32'd1));
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__f_reset_reqs$D_OUT )
                     begin  
                         RTL__near_mem__icache__v__h3949  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h3943  = RTL__near_mem__icache__v__h3949 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_reset && RTL__near_mem__icache__rg_cset_in_cache ==7'd127&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__f_reset_reqs$D_OUT )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_reset: Flushed", RTL__near_mem__icache__v__h3943 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_reset: Flushed", RTL__near_mem__icache__v__h3943 ,"I_MMU_Cache");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h4098  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h4092  = RTL__near_mem__icache__v__h4098 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL__near_mem__icache__v__h4092 ,"D_MMU_Cache", RTL__near_mem__icache__rg_addr );
                      else $display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL__near_mem__icache__v__h4092 ,"I_MMU_Cache", RTL__near_mem__icache__rg_addr );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        eaddr = {CTag 0x%0h  CSet 0x%0h  Word64 0x%0h  Byte 0x%0h}", RTL__near_mem__icache__pa_ctag__h4952 , RTL__near_mem__icache__rg_addr [11:5], RTL__near_mem__icache__rg_addr [4:3], RTL__near_mem__icache__rg_addr [2:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x: (state, tag):", RTL__near_mem__icache__rg_addr [11:5]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" (");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22])$write("CTAG_CLEAN");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22])$write("CTAG_EMPTY");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22])$write(", 0x%0x", RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [21:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22])$write(", --");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(")");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__icache__rg_addr [11:5], RTL__near_mem__icache__rg_addr [4:3]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" 0x%0x", RTL__near_mem__icache__ram_word64_set$DOB );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    TLB result: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_Xlate_Result { ","outcome: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_XLATE_OK");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","pa: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__rg_addr );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","exc_code: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'hA," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL__near_mem__icache__dmem_not_imem &&! RTL__near_mem__icache__soc_map$m_is_mem_addr && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => IO_REQ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$display("        Write-Cache-Hit: pa 0x%0h word64 0x%0h", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_st_amo_val );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        New Word64_Set:");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__icache__rg_addr [11:5], RTL__near_mem__icache__rg_addr [4:3]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write(" 0x%0x", RTL__near_mem__icache__IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op &&(! RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]||! RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Miss: pa 0x%0h word64 0x%0h", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_st_amo_val );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Hit/Miss: eaddr 0x%0h word64 0x%0h", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_st_amo_val );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__rg_op && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        => rl_write_response");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     begin  
                         RTL__near_mem__icache__v__h12540  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h12534  = RTL__near_mem__icache__v__h12540 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL__near_mem__icache__v__h12534 ,"D_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__word64__h5094 ,64'd0);
                      else $display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL__near_mem__icache__v__h12534 ,"I_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__word64__h5094 ,64'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&& RTL__near_mem__icache__NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )$display("        Read-hit: addr 0x%0h word64 0x%0h", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__word64__h5094 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL__near_mem__icache__dmem_not_imem || RTL__near_mem__icache__soc_map$m_is_mem_addr )&&! RTL__near_mem__icache__rg_op &&(! RTL__near_mem__icache__ram_state_and_ctag_cset$DOB [22]||! RTL__near_mem__icache__ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Read Miss: -> CACHE_START_REFILL.");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h14531  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h14525  = RTL__near_mem__icache__v__h14531 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_start_cache_refill: ", RTL__near_mem__icache__v__h14525 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_cache_refill: ", RTL__near_mem__icache__v__h14525 ,"I_MMU_Cache");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    To fabric: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__cline_fabric_addr__h14584 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd3);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'b011);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_cache_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    Victim way %0d; => CACHE_REFILL",1'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     begin  
                         RTL__near_mem__icache__v__h15336  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h15330  = RTL__near_mem__icache__v__h15336 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop:", RTL__near_mem__icache__v__h15330 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_cache_refill_rsps_loop:", RTL__near_mem__icache__v__h15330 ,"I_MMU_Cache");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rdata: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rresp: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rlast: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 &&! RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","ruser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h",1'd0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h15578  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h15572  = RTL__near_mem__icache__v__h15578 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL__near_mem__icache__v__h15572 ,"D_MMU_Cache", RTL__near_mem__icache__access_exc_code__h2256 );
                      else $display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL__near_mem__icache__v__h15572 ,"I_MMU_Cache", RTL__near_mem__icache__access_exc_code__h2256 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]==2'd3&&( RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL__near_mem__icache__rg_error_during_refill )&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => MODULE_EXCEPTION_RSP");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__rg_word64_set_in_cache [1:0]==2'd3&& RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0&&! RTL__near_mem__icache__rg_error_during_refill && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => CACHE_REREQ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$display("        Updating Cache word64_set 0x%0h, word64_in_cline %0d) old => new", RTL__near_mem__icache__rg_word64_set_in_cache , RTL__near_mem__icache__rg_word64_set_in_cache [1:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__icache__rg_addr [11:5], RTL__near_mem__icache__rg_word64_set_in_cache [1:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL__near_mem__icache__ram_word64_set$DOB );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL__near_mem__icache__rg_addr [11:5], RTL__near_mem__icache__rg_word64_set_in_cache [1:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_rereq && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL__near_mem__icache__rg_addr [11:5], RTL__near_mem__icache__rg_addr [11:3]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h17191  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h17185  = RTL__near_mem__icache__v__h17191 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL__near_mem__icache__v__h17185 ,"D_MMU_Cache", RTL__near_mem__icache__rg_f3 , RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_pa );
                      else $display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL__near_mem__icache__v__h17185 ,"I_MMU_Cache", RTL__near_mem__icache__rg_f3 , RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_pa );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__fabric_addr__h17243 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__value__h17372 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h17485  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h17479  = RTL__near_mem__icache__v__h17485 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL__near_mem__icache__v__h17479 ,"D_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_pa );
                      else $display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL__near_mem__icache__v__h17479 ,"I_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_pa );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rdata: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rresp: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rlast: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","ruser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h18585  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h18579  = RTL__near_mem__icache__v__h18585 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__icache__v__h18579 ,"D_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__ld_val__h17594 );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__icache__v__h18579 ,"I_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__ld_val__h17594 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h18692  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h18686  = RTL__near_mem__icache__v__h18692 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_read_rsp && RTL__near_mem__icache__master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL__near_mem__icache__v__h18686 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL__near_mem__icache__v__h18686 ,"I_MMU_Cache");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h18797  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h18791  = RTL__near_mem__icache__v__h18797 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__icache__v__h18791 ,"D_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_ld_val );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL__near_mem__icache__v__h18791 ,"I_MMU_Cache", RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_ld_val );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h18877  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h18871  = RTL__near_mem__icache__v__h18877 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL__near_mem__icache__v__h18871 ,"D_MMU_Cache", RTL__near_mem__icache__rg_f3 , RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_pa , RTL__near_mem__icache__rg_st_amo_val );
                      else $display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL__near_mem__icache__v__h18871 ,"I_MMU_Cache", RTL__near_mem__icache__rg_f3 , RTL__near_mem__icache__rg_addr , RTL__near_mem__icache__rg_pa , RTL__near_mem__icache__rg_st_amo_val );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_io_write_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => rl_ST_AMO_response");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h19505  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h19499  = RTL__near_mem__icache__v__h19505 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL__near_mem__icache__v__h19499 ,"D_MMU_Cache",$unsigned( RTL__near_mem__icache__b__h14485 ));
                      else $write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL__near_mem__icache__v__h19499 ,"I_MMU_Cache",$unsigned( RTL__near_mem__icache__b__h14485 ));
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","bresp: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","buser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     begin  
                         RTL__near_mem__icache__v__h19466  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h19460  = RTL__near_mem__icache__v__h19466 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL__near_mem__icache__v__h19460 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL__near_mem__icache__v__h19460 ,"I_MMU_Cache");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("    ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","bresp: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","buser: ");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h",1'd0," }");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_discard_write_rsp && RTL__near_mem__icache__master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h3483  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h3477  = RTL__near_mem__icache__v__h3483 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__WILL_FIRE_RL_rl_start_reset && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL__near_mem__icache__dmem_not_imem )$display("%0d: %s.rl_start_reset", RTL__near_mem__icache__v__h3477 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_reset", RTL__near_mem__icache__v__h3477 ,"I_MMU_Cache");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL__near_mem__icache__v__h19852  =$stime;#0;
                     end  
             RTL__near_mem__icache__v__h19846  = RTL__near_mem__icache__v__h19852 /32'd10;
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("%0d: %m.req: op:", RTL__near_mem__icache__v__h19846 );
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__req_op )$write("CACHE_ST");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL__near_mem__icache__req_op )$write("CACHE_LD");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" f3:%0d addr:0x%0h st_value:0x%0h", RTL__near_mem__icache__req_f3 , RTL__near_mem__icache__req_addr , RTL__near_mem__icache__req_st_value ,"\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    priv:");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__req_priv ==2'b0)$write("U");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__req_priv ==2'b01)$write("S");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__req_priv ==2'b11)$write("M");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL__near_mem__icache__req_priv !=2'b0&& RTL__near_mem__icache__req_priv !=2'b01&& RTL__near_mem__icache__req_priv !=2'b11)$write("RESERVED");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" sstatus_SUM:%0d mstatus_MXR:%0d satp:0x%0h", RTL__near_mem__icache__req_sstatus_SUM , RTL__near_mem__icache__req_mstatus_MXR , RTL__near_mem__icache__req_satp ,"\n");
             if ( RTL__near_mem__icache__RST_N !=1'b0)
                 if ( RTL__near_mem__icache__EN_req && RTL__near_mem__icache__req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 && RTL__near_mem__icache__NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL__near_mem__icache__req_addr [11:5], RTL__near_mem__icache__req_addr [11:3]);
         end
  assign  RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL__near_mem__icache__rg_addr ; 
  assign  RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL__near_mem__icache__rg_pa ;
    assign RTL__near_mem__CLK = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__RST_N = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache$mem_master_awready = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache$mem_master_bresp = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__dcache$mem_master_bvalid = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache$mem_master_rdata = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__dcache$mem_master_rid = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache$mem_master_rlast = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__dcache$mem_master_rresp = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache$mem_master_rvalid = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__dcache$mem_master_wready = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__dcache$req_addr = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__dcache$req_f3 = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__dcache$req_mstatus_MXR = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__dcache$EN_server_reset_response_get = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__dcache$valid = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL__near_mem__dcache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL__near_mem__dcache__CLK = RTL__near_mem__CLK;
    assign RTL__near_mem__dcache__RST_N = RTL__near_mem__RST_N;
    assign RTL__near_mem__dcache__set_verbosity_verbosity = RTL__near_mem__dcache$set_verbosity_verbosity;
    assign RTL__near_mem__dcache__EN_set_verbosity = RTL__near_mem__dcache$EN_set_verbosity;
    assign RTL__near_mem__dcache__EN_server_reset_request_put = RTL__near_mem__dcache$EN_server_reset_request_put;
    assign RTL__near_mem__dcache$RDY_server_reset_request_put = RTL__near_mem__dcache__RDY_server_reset_request_put;
    assign RTL__near_mem__dcache__EN_server_reset_response_get = RTL__near_mem__dcache$EN_server_reset_response_get;
    assign RTL__near_mem__dcache$RDY_server_reset_response_get = RTL__near_mem__dcache__RDY_server_reset_response_get;
    assign RTL__near_mem__dcache__req_op = RTL__near_mem__dcache$req_op;
    assign RTL__near_mem__dcache__req_f3 = RTL__near_mem__dcache$req_f3;
    assign RTL__near_mem__dcache__req_addr = RTL__near_mem__dcache$req_addr;
    assign RTL__near_mem__dcache__req_st_value = RTL__near_mem__dcache$req_st_value;
    assign RTL__near_mem__dcache__req_priv = RTL__near_mem__dcache$req_priv;
    assign RTL__near_mem__dcache__req_sstatus_SUM = RTL__near_mem__dcache$req_sstatus_SUM;
    assign RTL__near_mem__dcache__req_mstatus_MXR = RTL__near_mem__dcache$req_mstatus_MXR;
    assign RTL__near_mem__dcache__req_satp = RTL__near_mem__dcache$req_satp;
    assign RTL__near_mem__dcache__EN_req = RTL__near_mem__dcache$EN_req;
    assign RTL__near_mem__dcache$valid = RTL__near_mem__dcache__valid;
    assign RTL__near_mem__dcache$word64 = RTL__near_mem__dcache__word64;
    assign RTL__near_mem__dcache$exc = RTL__near_mem__dcache__exc;
    assign RTL__near_mem__dcache$exc_code = RTL__near_mem__dcache__exc_code;
    assign RTL__near_mem__dcache__EN_server_flush_request_put = RTL__near_mem__dcache$EN_server_flush_request_put;
    assign RTL__near_mem__dcache$RDY_server_flush_request_put = RTL__near_mem__dcache__RDY_server_flush_request_put;
    assign RTL__near_mem__dcache__EN_server_flush_response_get = RTL__near_mem__dcache$EN_server_flush_response_get;
    assign RTL__near_mem__dcache$RDY_server_flush_response_get = RTL__near_mem__dcache__RDY_server_flush_response_get;
    assign RTL__near_mem__dcache__EN_tlb_flush = RTL__near_mem__dcache$EN_tlb_flush;
    assign RTL__near_mem__dcache$mem_master_awvalid = RTL__near_mem__dcache__mem_master_awvalid;
    assign RTL__near_mem__dcache$mem_master_awid = RTL__near_mem__dcache__mem_master_awid;
    assign RTL__near_mem__dcache$mem_master_awaddr = RTL__near_mem__dcache__mem_master_awaddr;
    assign RTL__near_mem__dcache$mem_master_awlen = RTL__near_mem__dcache__mem_master_awlen;
    assign RTL__near_mem__dcache$mem_master_awsize = RTL__near_mem__dcache__mem_master_awsize;
    assign RTL__near_mem__dcache$mem_master_awburst = RTL__near_mem__dcache__mem_master_awburst;
    assign RTL__near_mem__dcache$mem_master_awlock = RTL__near_mem__dcache__mem_master_awlock;
    assign RTL__near_mem__dcache$mem_master_awcache = RTL__near_mem__dcache__mem_master_awcache;
    assign RTL__near_mem__dcache$mem_master_awprot = RTL__near_mem__dcache__mem_master_awprot;
    assign RTL__near_mem__dcache$mem_master_awqos = RTL__near_mem__dcache__mem_master_awqos;
    assign RTL__near_mem__dcache$mem_master_awregion = RTL__near_mem__dcache__mem_master_awregion;
    assign RTL__near_mem__dcache__mem_master_awready = RTL__near_mem__dcache$mem_master_awready;
    assign RTL__near_mem__dcache$mem_master_wvalid = RTL__near_mem__dcache__mem_master_wvalid;
    assign RTL__near_mem__dcache$mem_master_wdata = RTL__near_mem__dcache__mem_master_wdata;
    assign RTL__near_mem__dcache$mem_master_wstrb = RTL__near_mem__dcache__mem_master_wstrb;
    assign RTL__near_mem__dcache$mem_master_wlast = RTL__near_mem__dcache__mem_master_wlast;
    assign RTL__near_mem__dcache__mem_master_wready = RTL__near_mem__dcache$mem_master_wready;
    assign RTL__near_mem__dcache__mem_master_bvalid = RTL__near_mem__dcache$mem_master_bvalid;
    assign RTL__near_mem__dcache__mem_master_bid = RTL__near_mem__dcache$mem_master_bid;
    assign RTL__near_mem__dcache__mem_master_bresp = RTL__near_mem__dcache$mem_master_bresp;
    assign RTL__near_mem__dcache$mem_master_bready = RTL__near_mem__dcache__mem_master_bready;
    assign RTL__near_mem__dcache$mem_master_arvalid = RTL__near_mem__dcache__mem_master_arvalid;
    assign RTL__near_mem__icache$mem_master_arid = RTL__near_mem__icache__mem_master_arid;
    assign RTL__near_mem__icache$mem_master_araddr = RTL__near_mem__icache__mem_master_araddr;
    assign RTL__near_mem__icache$mem_master_arlen = RTL__near_mem__icache__mem_master_arlen;
    assign RTL__near_mem__icache$mem_master_arsize = RTL__near_mem__icache__mem_master_arsize;
    assign RTL__near_mem__icache$mem_master_arburst = RTL__near_mem__icache__mem_master_arburst;
    assign RTL__near_mem__icache$mem_master_arlock = RTL__near_mem__icache__mem_master_arlock;
    assign RTL__near_mem__icache$mem_master_arcache = RTL__near_mem__icache__mem_master_arcache;
    assign RTL__near_mem__icache$mem_master_arprot = RTL__near_mem__icache__mem_master_arprot;
    assign RTL__near_mem__icache$mem_master_arqos = RTL__near_mem__icache__mem_master_arqos;
    assign RTL__near_mem__icache$mem_master_arregion = RTL__near_mem__icache__mem_master_arregion;
    assign RTL__near_mem__icache__mem_master_arready = RTL__near_mem__icache$mem_master_arready;
    assign RTL__near_mem__icache__mem_master_rvalid = RTL__near_mem__icache$mem_master_rvalid;
    assign RTL__near_mem__icache__mem_master_rid = RTL__near_mem__icache$mem_master_rid;
    assign RTL__near_mem__icache__mem_master_rdata = RTL__near_mem__icache$mem_master_rdata;
    assign RTL__near_mem__icache__mem_master_rresp = RTL__near_mem__icache$mem_master_rresp;
    assign RTL__near_mem__icache__mem_master_rlast = RTL__near_mem__icache$mem_master_rlast;
    assign RTL__near_mem__icache$mem_master_rready = RTL__near_mem__icache__mem_master_rready;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache$req_satp = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__icache$req_st_value = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache$valid = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__near_mem__icache$addr = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__near_mem__icache$word64 = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache$exc = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__near_mem__icache$exc_code = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__near_mem__icache$RDY_server_flush_request_put = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__icache$RDY_server_flush_response_get = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__near_mem__icache$mem_master_awvalid = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache$mem_master_awid = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__near_mem__icache$mem_master_awaddr = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__near_mem__icache$mem_master_awlen = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__near_mem__icache$mem_master_awsize = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__near_mem__icache$mem_master_awburst = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL__near_mem__icache$mem_master_awlock = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__near_mem__icache$mem_master_awprot = RTL__near_mem__icache__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL__near_mem__icache__CLK = RTL__near_mem__CLK;
    assign RTL__near_mem__icache__RST_N = RTL__near_mem__RST_N;
    assign RTL__near_mem__icache__set_verbosity_verbosity = RTL__near_mem__icache$set_verbosity_verbosity;
    assign RTL__near_mem__icache__EN_set_verbosity = RTL__near_mem__icache$EN_set_verbosity;
    assign RTL__near_mem__icache__EN_server_reset_request_put = RTL__near_mem__icache$EN_server_reset_request_put;
    assign RTL__near_mem__icache$RDY_server_reset_request_put = RTL__near_mem__icache__RDY_server_reset_request_put;
    assign RTL__near_mem__icache__EN_server_reset_response_get = RTL__near_mem__icache$EN_server_reset_response_get;
    assign RTL__near_mem__icache$RDY_server_reset_response_get = RTL__near_mem__icache__RDY_server_reset_response_get;
    assign RTL__near_mem__icache__req_op = RTL__near_mem__icache$req_op;
    assign RTL__near_mem__icache__req_f3 = RTL__near_mem__icache$req_f3;
    assign RTL__near_mem__icache__req_addr = RTL__near_mem__icache$req_addr;
    assign RTL__near_mem__icache__req_st_value = RTL__near_mem__icache$req_st_value;
    assign RTL__near_mem__icache__req_priv = RTL__near_mem__icache$req_priv;
    assign RTL__near_mem__icache__req_sstatus_SUM = RTL__near_mem__icache$req_sstatus_SUM;
    assign RTL__near_mem__icache__req_mstatus_MXR = RTL__near_mem__icache$req_mstatus_MXR;
    assign RTL__near_mem__icache__req_satp = RTL__near_mem__icache$req_satp;
    assign RTL__near_mem__icache__EN_req = RTL__near_mem__icache$EN_req;
    assign RTL__near_mem__icache$valid = RTL__near_mem__icache__valid;
    assign RTL__near_mem__icache$addr = RTL__near_mem__icache__addr;
    assign RTL__near_mem__icache$word64 = RTL__near_mem__icache__word64;
    assign RTL__near_mem__icache$exc = RTL__near_mem__icache__exc;
    assign RTL__near_mem__icache$exc_code = RTL__near_mem__icache__exc_code;
    assign RTL__near_mem__icache__EN_server_flush_request_put = RTL__near_mem__icache$EN_server_flush_request_put;
    assign RTL__near_mem__icache$RDY_server_flush_request_put = RTL__near_mem__icache__RDY_server_flush_request_put;
    assign RTL__near_mem__icache__EN_server_flush_response_get = RTL__near_mem__icache$EN_server_flush_response_get;
    assign RTL__near_mem__icache$RDY_server_flush_response_get = RTL__near_mem__icache__RDY_server_flush_response_get;
    assign RTL__near_mem__icache__EN_tlb_flush = RTL__near_mem__icache$EN_tlb_flush;
    assign RTL__near_mem__icache$mem_master_awvalid = RTL__near_mem__icache__mem_master_awvalid;
    assign RTL__near_mem__icache$mem_master_awid = RTL__near_mem__icache__mem_master_awid;
    assign RTL__near_mem__icache$mem_master_awaddr = RTL__near_mem__icache__mem_master_awaddr;
    assign RTL__near_mem__icache$mem_master_awlen = RTL__near_mem__icache__mem_master_awlen;
    assign RTL__near_mem__icache$mem_master_awsize = RTL__near_mem__icache__mem_master_awsize;
      
    
    wire[63:0] RTL__near_mem__soc_map__m_boot_rom_addr_base , RTL__near_mem__soc_map__m_boot_rom_addr_lim , RTL__near_mem__soc_map__m_boot_rom_addr_size , RTL__near_mem__soc_map__m_mem0_controller_addr_base , RTL__near_mem__soc_map__m_mem0_controller_addr_lim , RTL__near_mem__soc_map__m_mem0_controller_addr_size , RTL__near_mem__soc_map__m_mtvec_reset_value , RTL__near_mem__soc_map__m_near_mem_io_addr_base , RTL__near_mem__soc_map__m_near_mem_io_addr_lim , RTL__near_mem__soc_map__m_near_mem_io_addr_size , RTL__near_mem__soc_map__m_nmivec_reset_value , RTL__near_mem__soc_map__m_pc_reset_value , RTL__near_mem__soc_map__m_plic_addr_base , RTL__near_mem__soc_map__m_plic_addr_lim , RTL__near_mem__soc_map__m_plic_addr_size , RTL__near_mem__soc_map__m_tcm_addr_base , RTL__near_mem__soc_map__m_tcm_addr_lim , RTL__near_mem__soc_map__m_tcm_addr_size , RTL__near_mem__soc_map__m_uart0_addr_base , RTL__near_mem__soc_map__m_uart0_addr_lim , RTL__near_mem__soc_map__m_uart0_addr_size ; 
    wire RTL__near_mem__soc_map__m_is_IO_addr , RTL__near_mem__soc_map__m_is_mem_addr , RTL__near_mem__soc_map__m_is_near_mem_IO_addr ; 
  assign  RTL__near_mem__soc_map__m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL__near_mem__soc_map__m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL__near_mem__soc_map__m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL__near_mem__soc_map__m_plic_addr_base =64'h000000000C000000; 
  assign  RTL__near_mem__soc_map__m_plic_addr_size =64'h0000000000400000; 
  assign  RTL__near_mem__soc_map__m_plic_addr_lim =64'd205520896; 
  assign  RTL__near_mem__soc_map__m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL__near_mem__soc_map__m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL__near_mem__soc_map__m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL__near_mem__soc_map__m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL__near_mem__soc_map__m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL__near_mem__soc_map__m_boot_rom_addr_lim =64'd8192; 
  assign  RTL__near_mem__soc_map__m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL__near_mem__soc_map__m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL__near_mem__soc_map__m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL__near_mem__soc_map__m_tcm_addr_base =64'h0; 
  assign  RTL__near_mem__soc_map__m_tcm_addr_size =64'd0; 
  assign  RTL__near_mem__soc_map__m_tcm_addr_lim =64'd0; 
  assign  RTL__near_mem__soc_map__m_is_mem_addr = RTL__near_mem__soc_map__m_is_mem_addr_addr >=64'h0000000000001000&& RTL__near_mem__soc_map__m_is_mem_addr_addr <64'd8192|| RTL__near_mem__soc_map__m_is_mem_addr_addr >=64'h0000000080000000&& RTL__near_mem__soc_map__m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL__near_mem__soc_map__m_is_IO_addr = RTL__near_mem__soc_map__m_is_IO_addr_addr >=64'h0000000002000000&& RTL__near_mem__soc_map__m_is_IO_addr_addr <64'd33603584|| RTL__near_mem__soc_map__m_is_IO_addr_addr >=64'h000000000C000000&& RTL__near_mem__soc_map__m_is_IO_addr_addr <64'd205520896|| RTL__near_mem__soc_map__m_is_IO_addr_addr >=64'h00000000C0000000&& RTL__near_mem__soc_map__m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL__near_mem__soc_map__m_is_near_mem_IO_addr = RTL__near_mem__soc_map__m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL__near_mem__soc_map__m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL__near_mem__soc_map__m_pc_reset_value =64'h0000000000001000; 
  assign  RTL__near_mem__soc_map__m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL__near_mem__soc_map__m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
    assign RTL__near_mem__dcache__soc_map__CLK = RTL__near_mem__dcache__CLK;
    assign RTL__near_mem__dcache__soc_map__RST_N = RTL__near_mem__dcache__RST_N;
    assign RTL__near_mem__dcache__soc_map__m_is_mem_addr_addr = RTL__near_mem__dcache__soc_map$m_is_mem_addr_addr;
    assign RTL__near_mem__dcache__soc_map$m_is_mem_addr = RTL__near_mem__dcache__soc_map__m_is_mem_addr;
    assign RTL__near_mem__dcache__soc_map__m_is_IO_addr_addr = RTL__near_mem__dcache__soc_map$m_is_IO_addr_addr;
    assign RTL__near_mem__dcache__soc_map__m_is_near_mem_IO_addr_addr = RTL__near_mem__dcache__soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL__near_mem__icache__soc_map__CLK = RTL__near_mem__icache__CLK;
    assign RTL__near_mem__icache__soc_map__RST_N = RTL__near_mem__icache__RST_N;
    assign RTL__near_mem__icache__soc_map__m_is_mem_addr_addr = RTL__near_mem__icache__soc_map$m_is_mem_addr_addr;
    assign RTL__near_mem__icache__soc_map$m_is_mem_addr = RTL__near_mem__icache__soc_map__m_is_mem_addr;
    assign RTL__near_mem__icache__soc_map__m_is_IO_addr_addr = RTL__near_mem__icache__soc_map$m_is_IO_addr_addr;
    assign RTL__near_mem__icache__soc_map__m_is_near_mem_IO_addr_addr = RTL__near_mem__icache__soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL__near_mem__soc_map__CLK = RTL__near_mem__CLK;
    assign RTL__near_mem__soc_map__RST_N = RTL__near_mem__RST_N;
    assign RTL__near_mem__soc_map__m_is_mem_addr_addr = RTL__near_mem__soc_map$m_is_mem_addr_addr;
    assign RTL__near_mem__soc_map__m_is_IO_addr_addr = RTL__near_mem__soc_map$m_is_IO_addr_addr;
    assign RTL__near_mem__soc_map__m_is_near_mem_IO_addr_addr = RTL__near_mem__soc_map$m_is_near_mem_IO_addr_addr;
     
  assign  RTL__near_mem__CAN_FIRE_RL_rl_reset = RTL__near_mem__dcache$RDY_server_reset_request_put && RTL__near_mem__icache$RDY_server_reset_request_put && RTL__near_mem__rg_state ==2'd0; 
  assign  RTL__near_mem__WILL_FIRE_RL_rl_reset = RTL__near_mem__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__CAN_FIRE_RL_rl_reset_complete = RTL__near_mem__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__WILL_FIRE_RL_rl_reset_complete = RTL__near_mem__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__MUX_rg_state$write_1__SEL_2 = RTL__near_mem__CAN_FIRE_RL_rl_reset &&! RTL__near_mem__EN_server_fence_request_put &&! RTL__near_mem__EN_server_fence_i_request_put ; 
  assign  RTL__near_mem__MUX_rg_state$write_1__SEL_3 = RTL__near_mem__dcache$RDY_server_reset_response_get && RTL__near_mem__icache$RDY_server_reset_response_get && RTL__near_mem__f_reset_rsps$FULL_N && RTL__near_mem__rg_state ==2'd1; 
  assign  RTL__near_mem__cfg_verbosity$D_IN =4'h0; 
  assign  RTL__near_mem__cfg_verbosity$EN =1'b0; 
  always @(    RTL__near_mem__EN_server_reset_request_put              or   RTL__near_mem__WILL_FIRE_RL_rl_reset           or   RTL__near_mem__WILL_FIRE_RL_rl_reset_complete  )
         begin 
             case (1'b1) 
              RTL__near_mem__EN_server_reset_request_put  : 
                  RTL__near_mem__rg_state$D_IN  =2'd0; 
              RTL__near_mem__WILL_FIRE_RL_rl_reset  : 
                  RTL__near_mem__rg_state$D_IN  =2'd1; 
              RTL__near_mem__WILL_FIRE_RL_rl_reset_complete  : 
                  RTL__near_mem__rg_state$D_IN  =2'd2;
              default : 
                  RTL__near_mem__rg_state$D_IN  =2'b10;endcase
         end
  assign  RTL__near_mem__rg_state$EN = RTL__near_mem__EN_server_reset_request_put || RTL__near_mem__WILL_FIRE_RL_rl_reset || RTL__near_mem__WILL_FIRE_RL_rl_reset_complete ; 
  assign  RTL__near_mem__dcache$mem_master_arready = RTL__near_mem__dmem_master_arready ; 
  assign  RTL__near_mem__dcache$mem_master_awready = RTL__near_mem__dmem_master_awready ; 
  assign  RTL__near_mem__dcache$mem_master_bid = RTL__near_mem__dmem_master_bid ; 
  assign  RTL__near_mem__dcache$mem_master_bresp = RTL__near_mem__dmem_master_bresp ; 
  assign  RTL__near_mem__dcache$mem_master_bvalid = RTL__near_mem__dmem_master_bvalid ; 
  assign  RTL__near_mem__dcache$mem_master_rdata = RTL__near_mem__dmem_master_rdata ; 
  assign  RTL__near_mem__dcache$mem_master_rid = RTL__near_mem__dmem_master_rid ; 
  assign  RTL__near_mem__dcache$mem_master_rlast = RTL__near_mem__dmem_master_rlast ; 
  assign  RTL__near_mem__dcache$mem_master_rresp = RTL__near_mem__dmem_master_rresp ; 
  assign  RTL__near_mem__dcache$mem_master_rvalid = RTL__near_mem__dmem_master_rvalid ; 
  assign  RTL__near_mem__dcache$mem_master_wready = RTL__near_mem__dmem_master_wready ; 
  assign  RTL__near_mem__dcache$req_addr = RTL__near_mem__dmem_req_addr ; 
  assign  RTL__near_mem__dcache$req_f3 = RTL__near_mem__dmem_req_f3 ; 
  assign  RTL__near_mem__dcache$req_mstatus_MXR = RTL__near_mem__dmem_req_mstatus_MXR ; 
  assign  RTL__near_mem__dcache$req_op = RTL__near_mem__dmem_req_op ; 
  assign  RTL__near_mem__dcache$req_priv = RTL__near_mem__dmem_req_priv ; 
  assign  RTL__near_mem__dcache$req_satp = RTL__near_mem__dmem_req_satp ; 
  assign  RTL__near_mem__dcache$req_sstatus_SUM = RTL__near_mem__dmem_req_sstatus_SUM ; 
  assign  RTL__near_mem__dcache$req_st_value = RTL__near_mem__dmem_req_store_value ; 
  assign  RTL__near_mem__dcache$set_verbosity_verbosity =4'h0; 
  assign  RTL__near_mem__dcache$EN_set_verbosity =1'b0; 
  assign  RTL__near_mem__dcache$EN_server_reset_request_put = RTL__near_mem__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__dcache$EN_server_reset_response_get = RTL__near_mem__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__dcache$EN_req = RTL__near_mem__EN_dmem_req ; 
  assign  RTL__near_mem__dcache$EN_server_flush_request_put = RTL__near_mem__EN_server_fence_i_request_put || RTL__near_mem__EN_server_fence_request_put ; 
  assign  RTL__near_mem__dcache$EN_server_flush_response_get = RTL__near_mem__EN_server_fence_i_response_get || RTL__near_mem__EN_server_fence_response_get ; 
  assign  RTL__near_mem__dcache$EN_tlb_flush = RTL__near_mem__EN_sfence_vma ; 
  assign  RTL__near_mem__f_reset_rsps$ENQ = RTL__near_mem__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__f_reset_rsps$DEQ = RTL__near_mem__EN_server_reset_response_get ; 
  assign  RTL__near_mem__f_reset_rsps$CLR =1'b0; 
  assign  RTL__near_mem__icache$mem_master_arready = RTL__near_mem__imem_master_arready ; 
  assign  RTL__near_mem__icache$mem_master_awready = RTL__near_mem__imem_master_awready ; 
  assign  RTL__near_mem__icache$mem_master_bid = RTL__near_mem__imem_master_bid ; 
  assign  RTL__near_mem__icache$mem_master_bresp = RTL__near_mem__imem_master_bresp ; 
  assign  RTL__near_mem__icache$mem_master_bvalid = RTL__near_mem__imem_master_bvalid ; 
  assign  RTL__near_mem__icache$mem_master_rdata = RTL__near_mem__imem_master_rdata ; 
  assign  RTL__near_mem__icache$mem_master_rid = RTL__near_mem__imem_master_rid ; 
  assign  RTL__near_mem__icache$mem_master_rlast = RTL__near_mem__imem_master_rlast ; 
  assign  RTL__near_mem__icache$mem_master_rresp = RTL__near_mem__imem_master_rresp ; 
  assign  RTL__near_mem__icache$mem_master_rvalid = RTL__near_mem__imem_master_rvalid ; 
  assign  RTL__near_mem__icache$mem_master_wready = RTL__near_mem__imem_master_wready ; 
  assign  RTL__near_mem__icache$req_addr = RTL__near_mem__imem_req_addr ; 
  assign  RTL__near_mem__icache$req_f3 = RTL__near_mem__imem_req_f3 ; 
  assign  RTL__near_mem__icache$req_mstatus_MXR = RTL__near_mem__imem_req_mstatus_MXR ; 
  assign  RTL__near_mem__icache$req_op =1'd0; 
  assign  RTL__near_mem__icache$req_priv = RTL__near_mem__imem_req_priv ; 
  assign  RTL__near_mem__icache$req_satp = RTL__near_mem__imem_req_satp ; 
  assign  RTL__near_mem__icache$req_sstatus_SUM = RTL__near_mem__imem_req_sstatus_SUM ; 
  assign  RTL__near_mem__icache$req_st_value =64'hAAAAAAAAAAAAAAAA; 
  assign  RTL__near_mem__icache$set_verbosity_verbosity =4'h0; 
  assign  RTL__near_mem__icache$EN_set_verbosity =1'b0; 
  assign  RTL__near_mem__icache$EN_server_reset_request_put = RTL__near_mem__MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL__near_mem__icache$EN_server_reset_response_get = RTL__near_mem__MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL__near_mem__icache$EN_req = RTL__near_mem__EN_imem_req ; 
  assign  RTL__near_mem__icache$EN_server_flush_request_put = RTL__near_mem__EN_server_fence_i_request_put ; 
  assign  RTL__near_mem__icache$EN_server_flush_response_get = RTL__near_mem__EN_server_fence_i_response_get ; 
  assign  RTL__near_mem__icache$EN_tlb_flush = RTL__near_mem__EN_sfence_vma ; 
  assign  RTL__near_mem__soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL__near_mem__soc_map$m_is_mem_addr_addr =64'h0; 
  assign  RTL__near_mem__soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL__near_mem__NOT_cfg_verbosity_read_ULE_1___d9 = RTL__near_mem__cfg_verbosity >4'd1; 
  always @( posedge  RTL__near_mem__CLK )
         begin 
             if ( RTL__near_mem__RST_N ==1'b0)
                 begin  
                     RTL__near_mem__cfg_verbosity  <=4'd0; 
                     RTL__near_mem__rg_state  <=2'd2;
                 end 
              else 
                 begin 
                     if ( RTL__near_mem__cfg_verbosity$EN ) 
                         RTL__near_mem__cfg_verbosity  <= RTL__near_mem__cfg_verbosity$D_IN ;
                     if ( RTL__near_mem__rg_state$EN ) 
                         RTL__near_mem__rg_state  <= RTL__near_mem__rg_state$D_IN ;
                 end 
         end
  always @( negedge  RTL__near_mem__CLK )
         begin #0;
             if ( RTL__near_mem__RST_N !=1'b0)
                 if ( RTL__near_mem__WILL_FIRE_RL_rl_reset && RTL__near_mem__NOT_cfg_verbosity_read_ULE_1___d9 )
                     begin  
                         RTL__near_mem__v__h1643  =$stime;#0;
                     end  
             RTL__near_mem__v__h1637  = RTL__near_mem__v__h1643 /32'd10;
             if ( RTL__near_mem__RST_N !=1'b0)
                 if ( RTL__near_mem__WILL_FIRE_RL_rl_reset && RTL__near_mem__NOT_cfg_verbosity_read_ULE_1___d9 )$display("%0d: Near_Mem.rl_reset", RTL__near_mem__v__h1637 );
             if ( RTL__near_mem__RST_N !=1'b0)
                 if ( RTL__near_mem__WILL_FIRE_RL_rl_reset_complete && RTL__near_mem__NOT_cfg_verbosity_read_ULE_1___d9 )
                     begin  
                         RTL__near_mem__v__h1794  =$stime;#0;
                     end  
             RTL__near_mem__v__h1788  = RTL__near_mem__v__h1794 /32'd10;
             if ( RTL__near_mem__RST_N !=1'b0)
                 if ( RTL__near_mem__WILL_FIRE_RL_rl_reset_complete && RTL__near_mem__NOT_cfg_verbosity_read_ULE_1___d9 )$display("%0d: Near_Mem.rl_reset_complete", RTL__near_mem__v__h1788 );
         end
 
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL__near_mem__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__near_mem__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__near_mem__CLK = RTL__CLK;
    assign RTL__near_mem__RST_N = RTL__RST_N;
    assign RTL__near_mem__EN_server_reset_request_put = RTL__near_mem$EN_server_reset_request_put;
    assign RTL__near_mem$RDY_server_reset_request_put = RTL__near_mem__RDY_server_reset_request_put;
    assign RTL__near_mem__EN_server_reset_response_get = RTL__near_mem$EN_server_reset_response_get;
    assign RTL__near_mem$RDY_server_reset_response_get = RTL__near_mem__RDY_server_reset_response_get;
    assign RTL__near_mem__imem_req_f3 = RTL__near_mem$imem_req_f3;
    assign RTL__near_mem__imem_req_addr = RTL__near_mem$imem_req_addr;
    assign RTL__near_mem__imem_req_priv = RTL__near_mem$imem_req_priv;
    assign RTL__near_mem__imem_req_sstatus_SUM = RTL__near_mem$imem_req_sstatus_SUM;
    assign RTL__near_mem__imem_req_mstatus_MXR = RTL__near_mem$imem_req_mstatus_MXR;
    assign RTL__near_mem__imem_req_satp = RTL__near_mem$imem_req_satp;
    assign RTL__near_mem__EN_imem_req = RTL__near_mem$EN_imem_req;
    assign RTL__near_mem$imem_valid = RTL__near_mem__imem_valid;
    assign RTL__near_mem$imem_is_i32_not_i16 = RTL__near_mem__imem_is_i32_not_i16;
    assign RTL__near_mem$imem_pc = RTL__near_mem__imem_pc;
    assign RTL__near_mem$imem_instr = RTL__near_mem__imem_instr;
    assign RTL__near_mem$imem_exc = RTL__near_mem__imem_exc;
    assign RTL__near_mem$imem_exc_code = RTL__near_mem__imem_exc_code;
    assign RTL__near_mem$imem_tval = RTL__near_mem__imem_tval;
    assign RTL__near_mem$imem_master_awvalid = RTL__near_mem__imem_master_awvalid;
    assign RTL__near_mem$imem_master_awid = RTL__near_mem__imem_master_awid;
    assign RTL__near_mem$imem_master_awaddr = RTL__near_mem__imem_master_awaddr;
    assign RTL__near_mem$imem_master_awlen = RTL__near_mem__imem_master_awlen;
    assign RTL__near_mem$imem_master_awsize = RTL__near_mem__imem_master_awsize;
    assign RTL__near_mem$imem_master_awburst = RTL__near_mem__imem_master_awburst;
    assign RTL__near_mem$imem_master_awlock = RTL__near_mem__imem_master_awlock;
    assign RTL__near_mem$imem_master_awcache = RTL__near_mem__imem_master_awcache;
    assign RTL__near_mem$imem_master_awprot = RTL__near_mem__imem_master_awprot;
    assign RTL__near_mem$imem_master_awqos = RTL__near_mem__imem_master_awqos;
    assign RTL__near_mem$imem_master_awregion = RTL__near_mem__imem_master_awregion;
    assign RTL__near_mem__imem_master_awready = RTL__near_mem$imem_master_awready;
    assign RTL__near_mem$imem_master_wvalid = RTL__near_mem__imem_master_wvalid;
    assign RTL__near_mem$imem_master_wdata = RTL__near_mem__imem_master_wdata;
    assign RTL__near_mem$imem_master_wstrb = RTL__near_mem__imem_master_wstrb;
    assign RTL__near_mem$imem_master_wlast = RTL__near_mem__imem_master_wlast;
    assign RTL__near_mem__imem_master_wready = RTL__near_mem$imem_master_wready;
    assign RTL__near_mem__imem_master_bvalid = RTL__near_mem$imem_master_bvalid;
    assign RTL__near_mem__imem_master_bid = RTL__near_mem$imem_master_bid;
    assign RTL__near_mem__imem_master_bresp = RTL__near_mem$imem_master_bresp;
    assign RTL__near_mem$imem_master_bready = RTL__near_mem__imem_master_bready;
    assign RTL__near_mem$imem_master_arvalid = RTL__near_mem__imem_master_arvalid;
    assign RTL__near_mem$imem_master_arid = RTL__near_mem__imem_master_arid;
    assign RTL__near_mem$imem_master_araddr = RTL__near_mem__imem_master_araddr;
    assign RTL__near_mem$imem_master_arlen = RTL__near_mem__imem_master_arlen;
    assign RTL__near_mem$imem_master_arsize = RTL__near_mem__imem_master_arsize;
    assign RTL__near_mem$imem_master_arburst = RTL__near_mem__imem_master_arburst;
    assign RTL__near_mem$imem_master_arlock = RTL__near_mem__imem_master_arlock;
    assign RTL__near_mem$imem_master_arcache = RTL__near_mem__imem_master_arcache;
    assign RTL__near_mem$imem_master_arprot = RTL__near_mem__imem_master_arprot;
    assign RTL__near_mem$imem_master_arqos = RTL__near_mem__imem_master_arqos;
    assign RTL__near_mem$imem_master_arregion = RTL__near_mem__imem_master_arregion;
    assign RTL__near_mem__imem_master_arready = RTL__near_mem$imem_master_arready;
    assign RTL__near_mem__imem_master_rvalid = RTL__near_mem$imem_master_rvalid;
    assign RTL__near_mem__imem_master_rid = RTL__near_mem$imem_master_rid;
    assign RTL__near_mem__imem_master_rdata = RTL__near_mem$imem_master_rdata;
    assign RTL__near_mem__imem_master_rresp = RTL__near_mem$imem_master_rresp;
    assign RTL__near_mem__imem_master_rlast = RTL__near_mem$imem_master_rlast;
    assign RTL__near_mem$imem_master_rready = RTL__near_mem__imem_master_rready;
    assign RTL__near_mem__dmem_req_op = RTL__near_mem$dmem_req_op;
    assign RTL__near_mem__dmem_req_f3 = RTL__near_mem$dmem_req_f3;
    assign RTL__near_mem__dmem_req_addr = RTL__near_mem$dmem_req_addr;
    assign RTL__near_mem__dmem_req_store_value = RTL__near_mem$dmem_req_store_value;
    assign RTL__near_mem__dmem_req_priv = RTL__near_mem$dmem_req_priv;
    assign RTL__near_mem__dmem_req_sstatus_SUM = RTL__near_mem$dmem_req_sstatus_SUM;
    assign RTL__near_mem__dmem_req_mstatus_MXR = RTL__near_mem$dmem_req_mstatus_MXR;
    assign RTL__near_mem__dmem_req_satp = RTL__near_mem$dmem_req_satp;
    assign RTL__near_mem__EN_dmem_req = RTL__near_mem$EN_dmem_req;
    assign RTL__near_mem$dmem_valid = RTL__near_mem__dmem_valid;
    assign RTL__near_mem$dmem_word64 = RTL__near_mem__dmem_word64;
    assign RTL__near_mem$dmem_exc = RTL__near_mem__dmem_exc;
    assign RTL__near_mem$dmem_exc_code = RTL__near_mem__dmem_exc_code;
    assign RTL__near_mem$dmem_master_awvalid = RTL__near_mem__dmem_master_awvalid;
    assign RTL__near_mem$dmem_master_awid = RTL__near_mem__dmem_master_awid;
    assign RTL__near_mem$dmem_master_awaddr = RTL__near_mem__dmem_master_awaddr;
    assign RTL__near_mem$dmem_master_awlen = RTL__near_mem__dmem_master_awlen;
    assign RTL__near_mem$dmem_master_awsize = RTL__near_mem__dmem_master_awsize;
    assign RTL__near_mem$dmem_master_awburst = RTL__near_mem__dmem_master_awburst;
    assign RTL__near_mem$dmem_master_awlock = RTL__near_mem__dmem_master_awlock;
    assign RTL__near_mem$dmem_master_awcache = RTL__near_mem__dmem_master_awcache;
    assign RTL__near_mem$dmem_master_awprot = RTL__near_mem__dmem_master_awprot;
    assign RTL__near_mem$dmem_master_awqos = RTL__near_mem__dmem_master_awqos;
    assign RTL__near_mem$dmem_master_awregion = RTL__near_mem__dmem_master_awregion;
    assign RTL__near_mem__dmem_master_awready = RTL__near_mem$dmem_master_awready;
    assign RTL__near_mem$dmem_master_wvalid = RTL__near_mem__dmem_master_wvalid;
    assign RTL__near_mem$dmem_master_wdata = RTL__near_mem__dmem_master_wdata;
    assign RTL__near_mem$dmem_master_wstrb = RTL__near_mem__dmem_master_wstrb;
    assign RTL__near_mem$dmem_master_wlast = RTL__near_mem__dmem_master_wlast;
    assign RTL__near_mem__dmem_master_wready = RTL__near_mem$dmem_master_wready;
    assign RTL__near_mem__dmem_master_bvalid = RTL__near_mem$dmem_master_bvalid;
    assign RTL__near_mem__dmem_master_bid = RTL__near_mem$dmem_master_bid;
    assign RTL__near_mem__dmem_master_bresp = RTL__near_mem$dmem_master_bresp;
    assign RTL__near_mem$dmem_master_bready = RTL__near_mem__dmem_master_bready;
    assign RTL__near_mem$dmem_master_arvalid = RTL__near_mem__dmem_master_arvalid;
    assign RTL__near_mem$dmem_master_arid = RTL__near_mem__dmem_master_arid;
    assign RTL__near_mem$dmem_master_araddr = RTL__near_mem__dmem_master_araddr;
    assign RTL__near_mem$dmem_master_arlen = RTL__near_mem__dmem_master_arlen;
    assign RTL__near_mem$dmem_master_arsize = RTL__near_mem__dmem_master_arsize;
    assign RTL__near_mem$dmem_master_arburst = RTL__near_mem__dmem_master_arburst;
    assign RTL__near_mem$dmem_master_arlock = RTL__near_mem__dmem_master_arlock;
    assign RTL__near_mem$dmem_master_arcache = RTL__near_mem__dmem_master_arcache;
    assign RTL__near_mem$dmem_master_arprot = RTL__near_mem__dmem_master_arprot;
    assign RTL__near_mem$dmem_master_arqos = RTL__near_mem__dmem_master_arqos;
    assign RTL__near_mem$dmem_master_arregion = RTL__near_mem__dmem_master_arregion;
    assign RTL__near_mem__dmem_master_arready = RTL__near_mem$dmem_master_arready;
    assign RTL__near_mem__dmem_master_rvalid = RTL__near_mem$dmem_master_rvalid;
    assign RTL__near_mem__dmem_master_rid = RTL__near_mem$dmem_master_rid;
    assign RTL__near_mem__dmem_master_rdata = RTL__near_mem$dmem_master_rdata;
    assign RTL__near_mem__dmem_master_rresp = RTL__near_mem$dmem_master_rresp;
    assign RTL__near_mem__dmem_master_rlast = RTL__near_mem$dmem_master_rlast;
    assign RTL__near_mem$dmem_master_rready = RTL__near_mem__dmem_master_rready;
    assign RTL__near_mem__EN_server_fence_i_request_put = RTL__near_mem$EN_server_fence_i_request_put;
    assign RTL__near_mem$RDY_server_fence_i_request_put = RTL__near_mem__RDY_server_fence_i_request_put;
    assign RTL__near_mem__EN_server_fence_i_response_get = RTL__near_mem$EN_server_fence_i_response_get;
    assign RTL__near_mem$RDY_server_fence_i_response_get = RTL__near_mem__RDY_server_fence_i_response_get;
    assign RTL__near_mem__server_fence_request_put = RTL__near_mem$server_fence_request_put;
    assign RTL__near_mem__EN_server_fence_request_put = RTL__near_mem$EN_server_fence_request_put;
    assign RTL__near_mem$RDY_server_fence_request_put = RTL__near_mem__RDY_server_fence_request_put;
    assign RTL__near_mem__EN_server_fence_response_get = RTL__near_mem$EN_server_fence_response_get;
    assign RTL__near_mem$RDY_server_fence_response_get = RTL__near_mem__RDY_server_fence_response_get;
    assign RTL__near_mem__EN_sfence_vma = RTL__near_mem$EN_sfence_vma;
      
    
    wire[63:0] RTL__soc_map__m_boot_rom_addr_base , RTL__soc_map__m_boot_rom_addr_lim , RTL__soc_map__m_boot_rom_addr_size , RTL__soc_map__m_mem0_controller_addr_base , RTL__soc_map__m_mem0_controller_addr_lim , RTL__soc_map__m_mem0_controller_addr_size , RTL__soc_map__m_mtvec_reset_value , RTL__soc_map__m_near_mem_io_addr_base , RTL__soc_map__m_near_mem_io_addr_lim , RTL__soc_map__m_near_mem_io_addr_size , RTL__soc_map__m_nmivec_reset_value , RTL__soc_map__m_pc_reset_value , RTL__soc_map__m_plic_addr_base , RTL__soc_map__m_plic_addr_lim , RTL__soc_map__m_plic_addr_size , RTL__soc_map__m_tcm_addr_base , RTL__soc_map__m_tcm_addr_lim , RTL__soc_map__m_tcm_addr_size , RTL__soc_map__m_uart0_addr_base , RTL__soc_map__m_uart0_addr_lim , RTL__soc_map__m_uart0_addr_size ; 
    wire RTL__soc_map__m_is_IO_addr , RTL__soc_map__m_is_mem_addr , RTL__soc_map__m_is_near_mem_IO_addr ; 
  assign  RTL__soc_map__m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL__soc_map__m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL__soc_map__m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL__soc_map__m_plic_addr_base =64'h000000000C000000; 
  assign  RTL__soc_map__m_plic_addr_size =64'h0000000000400000; 
  assign  RTL__soc_map__m_plic_addr_lim =64'd205520896; 
  assign  RTL__soc_map__m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL__soc_map__m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL__soc_map__m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL__soc_map__m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL__soc_map__m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL__soc_map__m_boot_rom_addr_lim =64'd8192; 
  assign  RTL__soc_map__m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL__soc_map__m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL__soc_map__m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL__soc_map__m_tcm_addr_base =64'h0; 
  assign  RTL__soc_map__m_tcm_addr_size =64'd0; 
  assign  RTL__soc_map__m_tcm_addr_lim =64'd0; 
  assign  RTL__soc_map__m_is_mem_addr = RTL__soc_map__m_is_mem_addr_addr >=64'h0000000000001000&& RTL__soc_map__m_is_mem_addr_addr <64'd8192|| RTL__soc_map__m_is_mem_addr_addr >=64'h0000000080000000&& RTL__soc_map__m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL__soc_map__m_is_IO_addr = RTL__soc_map__m_is_IO_addr_addr >=64'h0000000002000000&& RTL__soc_map__m_is_IO_addr_addr <64'd33603584|| RTL__soc_map__m_is_IO_addr_addr >=64'h000000000C000000&& RTL__soc_map__m_is_IO_addr_addr <64'd205520896|| RTL__soc_map__m_is_IO_addr_addr >=64'h00000000C0000000&& RTL__soc_map__m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL__soc_map__m_is_near_mem_IO_addr = RTL__soc_map__m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL__soc_map__m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL__soc_map__m_pc_reset_value =64'h0000000000001000; 
  assign  RTL__soc_map__m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL__soc_map__m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
    assign RTL__csr_regfile__soc_map__CLK = RTL__csr_regfile__CLK;
    assign RTL__csr_regfile__soc_map__RST_N = RTL__csr_regfile__RST_N;
    assign RTL__csr_regfile__soc_map__m_is_mem_addr_addr = RTL__csr_regfile__soc_map$m_is_mem_addr_addr;
    assign RTL__csr_regfile__soc_map__m_is_IO_addr_addr = RTL__csr_regfile__soc_map$m_is_IO_addr_addr;
    assign RTL__csr_regfile__soc_map__m_is_near_mem_IO_addr_addr = RTL__csr_regfile__soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL__csr_regfile__soc_map$m_mtvec_reset_value = RTL__csr_regfile__soc_map__m_mtvec_reset_value;
    assign RTL__csr_regfile__soc_map$m_nmivec_reset_value = RTL__csr_regfile__soc_map__m_nmivec_reset_value;
    assign RTL__soc_map__CLK = RTL__CLK;
    assign RTL__soc_map__RST_N = RTL__RST_N;
    assign RTL__soc_map__m_is_mem_addr_addr = RTL__soc_map$m_is_mem_addr_addr;
    assign RTL__soc_map__m_is_IO_addr_addr = RTL__soc_map$m_is_IO_addr_addr;
    assign RTL__soc_map__m_is_near_mem_IO_addr_addr = RTL__soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL__soc_map$m_pc_reset_value = RTL__soc_map__m_pc_reset_value;
      
    
    parameter RTL__stage1_f_reset_reqs__guarded =1; 
    reg RTL__stage1_f_reset_reqs__empty_reg ; 
    reg RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__FULL_N = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__EMPTY_N = RTL__stage1_f_reset_reqs__empty_reg ; 
  always @( posedge  RTL__stage1_f_reset_reqs__CLK )
         begin 
             if ( RTL__stage1_f_reset_reqs__RST ==1'b0)
                 begin  
                     RTL__stage1_f_reset_reqs__empty_reg  <=1'b0; 
                     RTL__stage1_f_reset_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__stage1_f_reset_reqs__CLR )
                         begin  
                             RTL__stage1_f_reset_reqs__empty_reg  <=1'b0; 
                             RTL__stage1_f_reset_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__stage1_f_reset_reqs__ENQ &&! RTL__stage1_f_reset_reqs__DEQ )
                             begin  
                                 RTL__stage1_f_reset_reqs__empty_reg  <=1'b1; 
                                 RTL__stage1_f_reset_reqs__full_reg  <=! RTL__stage1_f_reset_reqs__empty_reg ;
                             end 
                          else 
                             if (! RTL__stage1_f_reset_reqs__ENQ && RTL__stage1_f_reset_reqs__DEQ )
                                 begin  
                                     RTL__stage1_f_reset_reqs__full_reg  <=1'b1; 
                                     RTL__stage1_f_reset_reqs__empty_reg  <=! RTL__stage1_f_reset_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__stage1_f_reset_reqs__CLK )
         begin : RTL__stage1_f_reset_reqs__error_checks 
           reg RTL__stage1_f_reset_reqs__deqerror , RTL__stage1_f_reset_reqs__enqerror ; 
             RTL__stage1_f_reset_reqs__deqerror  =0; 
             RTL__stage1_f_reset_reqs__enqerror  =0;
             if ( RTL__stage1_f_reset_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__stage1_f_reset_reqs__empty_reg && RTL__stage1_f_reset_reqs__DEQ )
                         begin  
                             RTL__stage1_f_reset_reqs__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__stage1_f_reset_reqs__full_reg && RTL__stage1_f_reset_reqs__ENQ &&(! RTL__stage1_f_reset_reqs__DEQ || RTL__stage1_f_reset_reqs__guarded ))
                         begin  
                             RTL__stage1_f_reset_reqs__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_reqs__full_reg ; 
  assign  RTL__stage1_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_reqs__empty_reg ;
    parameter RTL__stage1_f_reset_rsps__guarded =1; 
    reg RTL__stage1_f_reset_rsps__empty_reg ; 
    reg RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__FULL_N = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__EMPTY_N = RTL__stage1_f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__stage1_f_reset_rsps__CLK )
         begin 
             if ( RTL__stage1_f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__stage1_f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__stage1_f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__stage1_f_reset_rsps__CLR )
                         begin  
                             RTL__stage1_f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__stage1_f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__stage1_f_reset_rsps__ENQ &&! RTL__stage1_f_reset_rsps__DEQ )
                             begin  
                                 RTL__stage1_f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__stage1_f_reset_rsps__full_reg  <=! RTL__stage1_f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if (! RTL__stage1_f_reset_rsps__ENQ && RTL__stage1_f_reset_rsps__DEQ )
                                 begin  
                                     RTL__stage1_f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__stage1_f_reset_rsps__empty_reg  <=! RTL__stage1_f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__stage1_f_reset_rsps__CLK )
         begin : RTL__stage1_f_reset_rsps__error_checks 
           reg RTL__stage1_f_reset_rsps__deqerror , RTL__stage1_f_reset_rsps__enqerror ; 
             RTL__stage1_f_reset_rsps__deqerror  =0; 
             RTL__stage1_f_reset_rsps__enqerror  =0;
             if ( RTL__stage1_f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__stage1_f_reset_rsps__empty_reg && RTL__stage1_f_reset_rsps__DEQ )
                         begin  
                             RTL__stage1_f_reset_rsps__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__stage1_f_reset_rsps__full_reg && RTL__stage1_f_reset_rsps__ENQ &&(! RTL__stage1_f_reset_rsps__DEQ || RTL__stage1_f_reset_rsps__guarded ))
                         begin  
                             RTL__stage1_f_reset_rsps__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__stage1_f_reset_rsps__full_reg ; 
  assign  RTL__stage1_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage1_f_reset_rsps__empty_reg ;
    parameter RTL__stage2_f_reset_reqs__guarded =1; 
    reg RTL__stage2_f_reset_reqs__empty_reg ; 
    reg RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__FULL_N = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__EMPTY_N = RTL__stage2_f_reset_reqs__empty_reg ; 
  always @( posedge  RTL__stage2_f_reset_reqs__CLK )
         begin 
             if ( RTL__stage2_f_reset_reqs__RST ==1'b0)
                 begin  
                     RTL__stage2_f_reset_reqs__empty_reg  <=1'b0; 
                     RTL__stage2_f_reset_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__stage2_f_reset_reqs__CLR )
                         begin  
                             RTL__stage2_f_reset_reqs__empty_reg  <=1'b0; 
                             RTL__stage2_f_reset_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__stage2_f_reset_reqs__ENQ &&! RTL__stage2_f_reset_reqs__DEQ )
                             begin  
                                 RTL__stage2_f_reset_reqs__empty_reg  <=1'b1; 
                                 RTL__stage2_f_reset_reqs__full_reg  <=! RTL__stage2_f_reset_reqs__empty_reg ;
                             end 
                          else 
                             if (! RTL__stage2_f_reset_reqs__ENQ && RTL__stage2_f_reset_reqs__DEQ )
                                 begin  
                                     RTL__stage2_f_reset_reqs__full_reg  <=1'b1; 
                                     RTL__stage2_f_reset_reqs__empty_reg  <=! RTL__stage2_f_reset_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__stage2_f_reset_reqs__CLK )
         begin : RTL__stage2_f_reset_reqs__error_checks 
           reg RTL__stage2_f_reset_reqs__deqerror , RTL__stage2_f_reset_reqs__enqerror ; 
             RTL__stage2_f_reset_reqs__deqerror  =0; 
             RTL__stage2_f_reset_reqs__enqerror  =0;
             if ( RTL__stage2_f_reset_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__stage2_f_reset_reqs__empty_reg && RTL__stage2_f_reset_reqs__DEQ )
                         begin  
                             RTL__stage2_f_reset_reqs__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__stage2_f_reset_reqs__full_reg && RTL__stage2_f_reset_reqs__ENQ &&(! RTL__stage2_f_reset_reqs__DEQ || RTL__stage2_f_reset_reqs__guarded ))
                         begin  
                             RTL__stage2_f_reset_reqs__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_reqs__full_reg ; 
  assign  RTL__stage2_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_reqs__empty_reg ;
    parameter RTL__stage2_f_reset_rsps__guarded =1; 
    reg RTL__stage2_f_reset_rsps__empty_reg ; 
    reg RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__FULL_N = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__EMPTY_N = RTL__stage2_f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__stage2_f_reset_rsps__CLK )
         begin 
             if ( RTL__stage2_f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__stage2_f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__stage2_f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__stage2_f_reset_rsps__CLR )
                         begin  
                             RTL__stage2_f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__stage2_f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__stage2_f_reset_rsps__ENQ &&! RTL__stage2_f_reset_rsps__DEQ )
                             begin  
                                 RTL__stage2_f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__stage2_f_reset_rsps__full_reg  <=! RTL__stage2_f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if (! RTL__stage2_f_reset_rsps__ENQ && RTL__stage2_f_reset_rsps__DEQ )
                                 begin  
                                     RTL__stage2_f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__stage2_f_reset_rsps__empty_reg  <=! RTL__stage2_f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__stage2_f_reset_rsps__CLK )
         begin : RTL__stage2_f_reset_rsps__error_checks 
           reg RTL__stage2_f_reset_rsps__deqerror , RTL__stage2_f_reset_rsps__enqerror ; 
             RTL__stage2_f_reset_rsps__deqerror  =0; 
             RTL__stage2_f_reset_rsps__enqerror  =0;
             if ( RTL__stage2_f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__stage2_f_reset_rsps__empty_reg && RTL__stage2_f_reset_rsps__DEQ )
                         begin  
                             RTL__stage2_f_reset_rsps__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__stage2_f_reset_rsps__full_reg && RTL__stage2_f_reset_rsps__ENQ &&(! RTL__stage2_f_reset_rsps__DEQ || RTL__stage2_f_reset_rsps__guarded ))
                         begin  
                             RTL__stage2_f_reset_rsps__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__full_reg ; 
  assign  RTL__stage2_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__empty_reg ;
    parameter RTL__stage3_f_reset_reqs__guarded =1; 
    reg RTL__stage3_f_reset_reqs__empty_reg ; 
    reg RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__FULL_N = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__EMPTY_N = RTL__stage3_f_reset_reqs__empty_reg ; 
  always @( posedge  RTL__stage3_f_reset_reqs__CLK )
         begin 
             if ( RTL__stage3_f_reset_reqs__RST ==1'b0)
                 begin  
                     RTL__stage3_f_reset_reqs__empty_reg  <=1'b0; 
                     RTL__stage3_f_reset_reqs__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__stage3_f_reset_reqs__CLR )
                         begin  
                             RTL__stage3_f_reset_reqs__empty_reg  <=1'b0; 
                             RTL__stage3_f_reset_reqs__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__stage3_f_reset_reqs__ENQ &&! RTL__stage3_f_reset_reqs__DEQ )
                             begin  
                                 RTL__stage3_f_reset_reqs__empty_reg  <=1'b1; 
                                 RTL__stage3_f_reset_reqs__full_reg  <=! RTL__stage3_f_reset_reqs__empty_reg ;
                             end 
                          else 
                             if (! RTL__stage3_f_reset_reqs__ENQ && RTL__stage3_f_reset_reqs__DEQ )
                                 begin  
                                     RTL__stage3_f_reset_reqs__full_reg  <=1'b1; 
                                     RTL__stage3_f_reset_reqs__empty_reg  <=! RTL__stage3_f_reset_reqs__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__stage3_f_reset_reqs__CLK )
         begin : RTL__stage3_f_reset_reqs__error_checks 
           reg RTL__stage3_f_reset_reqs__deqerror , RTL__stage3_f_reset_reqs__enqerror ; 
             RTL__stage3_f_reset_reqs__deqerror  =0; 
             RTL__stage3_f_reset_reqs__enqerror  =0;
             if ( RTL__stage3_f_reset_reqs__RST ==!1'b0)
                 begin 
                     if (! RTL__stage3_f_reset_reqs__empty_reg && RTL__stage3_f_reset_reqs__DEQ )
                         begin  
                             RTL__stage3_f_reset_reqs__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__stage3_f_reset_reqs__full_reg && RTL__stage3_f_reset_reqs__ENQ &&(! RTL__stage3_f_reset_reqs__DEQ || RTL__stage3_f_reset_reqs__guarded ))
                         begin  
                             RTL__stage3_f_reset_reqs__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_reqs__full_reg ; 
  assign  RTL__stage3_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_reqs__empty_reg ;
    parameter RTL__stage3_f_reset_rsps__guarded =1; 
    reg RTL__stage3_f_reset_rsps__empty_reg ; 
    reg RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__FULL_N = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__EMPTY_N = RTL__stage3_f_reset_rsps__empty_reg ; 
  always @( posedge  RTL__stage3_f_reset_rsps__CLK )
         begin 
             if ( RTL__stage3_f_reset_rsps__RST ==1'b0)
                 begin  
                     RTL__stage3_f_reset_rsps__empty_reg  <=1'b0; 
                     RTL__stage3_f_reset_rsps__full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL__stage3_f_reset_rsps__CLR )
                         begin  
                             RTL__stage3_f_reset_rsps__empty_reg  <=1'b0; 
                             RTL__stage3_f_reset_rsps__full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL__stage3_f_reset_rsps__ENQ &&! RTL__stage3_f_reset_rsps__DEQ )
                             begin  
                                 RTL__stage3_f_reset_rsps__empty_reg  <=1'b1; 
                                 RTL__stage3_f_reset_rsps__full_reg  <=! RTL__stage3_f_reset_rsps__empty_reg ;
                             end 
                          else 
                             if (! RTL__stage3_f_reset_rsps__ENQ && RTL__stage3_f_reset_rsps__DEQ )
                                 begin  
                                     RTL__stage3_f_reset_rsps__full_reg  <=1'b1; 
                                     RTL__stage3_f_reset_rsps__empty_reg  <=! RTL__stage3_f_reset_rsps__full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL__stage3_f_reset_rsps__CLK )
         begin : RTL__stage3_f_reset_rsps__error_checks 
           reg RTL__stage3_f_reset_rsps__deqerror , RTL__stage3_f_reset_rsps__enqerror ; 
             RTL__stage3_f_reset_rsps__deqerror  =0; 
             RTL__stage3_f_reset_rsps__enqerror  =0;
             if ( RTL__stage3_f_reset_rsps__RST ==!1'b0)
                 begin 
                     if (! RTL__stage3_f_reset_rsps__empty_reg && RTL__stage3_f_reset_rsps__DEQ )
                         begin  
                             RTL__stage3_f_reset_rsps__deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL__stage3_f_reset_rsps__full_reg && RTL__stage3_f_reset_rsps__ENQ &&(! RTL__stage3_f_reset_rsps__DEQ || RTL__stage3_f_reset_rsps__guarded ))
                         begin  
                             RTL__stage3_f_reset_rsps__enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__full_reg ; 
  assign  RTL__stage3_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__empty_reg ;
    assign RTL__csr_regfile__f_reset_rsps__RST = RTL__csr_regfile__RST_N;
    assign RTL__csr_regfile__f_reset_rsps__CLK = RTL__csr_regfile__CLK;
    assign RTL__csr_regfile__f_reset_rsps__ENQ = RTL__csr_regfile__f_reset_rsps$ENQ;
    assign RTL__csr_regfile__f_reset_rsps__CLR = RTL__csr_regfile__f_reset_rsps$CLR;
    assign RTL__csr_regfile__f_reset_rsps__DEQ = RTL__csr_regfile__f_reset_rsps$DEQ;
    assign RTL__csr_regfile__f_reset_rsps$FULL_N = RTL__csr_regfile__f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__csr_regfile__f_reset_rsps$EMPTY_N = RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__csr_regfile__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__csr_regfile__f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    assign RTL__CLK = RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    assign RTL__stage1_f_reset_reqs$ENQ = RTL__stage1_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__stage1_f_reset_reqs$DEQ = RTL__stage1_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__stage1_f_reset_reqs$CLR = RTL__stage1_f_reset_reqs__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    assign RTL__stage1_f_reset_reqs$FULL_N = RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    assign RTL__stage1_f_reset_reqs$EMPTY_N = RTL__stage1_f_reset_reqs__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__stage1_f_reset_reqs__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__stage1_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    assign RTL__RST_N = RTL__stage1_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__CLK = RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    assign RTL__stage1_f_reset_rsps$ENQ = RTL__stage1_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    assign RTL__stage1_f_reset_rsps$DEQ = RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    assign RTL__stage1_f_reset_rsps$CLR = RTL__stage1_f_reset_rsps__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    assign RTL__stage1_f_reset_rsps$FULL_N = RTL__stage1_f_reset_rsps__FULL_N;
    assign RTL__stage1_f_reset_rsps$EMPTY_N = RTL__stage1_f_reset_rsps__EMPTY_N;
    assign RTL__stage1_f_reset_rsps__RST = RTL__RST_N;
    assign RTL__stage1_f_reset_rsps__CLK = RTL__CLK;
    assign RTL__stage2_f_reset_reqs__ENQ = RTL__stage2_f_reset_reqs$ENQ;
    assign RTL__stage2_f_reset_reqs__CLR = RTL__stage2_f_reset_reqs$CLR;
    assign RTL__stage2_f_reset_reqs__DEQ = RTL__stage2_f_reset_reqs$DEQ;
    assign RTL__stage2_f_reset_reqs$DEQ = RTL__stage2_f_reset_reqs__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__stage2_f_reset_reqs$CLR = RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__stage2_f_reset_reqs$FULL_N = RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__stage2_f_reset_reqs$EMPTY_N = RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__stage2_f_reset_reqs__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    assign RTL__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__stage2_f_reset_reqs__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    assign RTL__RST_N = RTL__stage2_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__CLK = RTL__stage2_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__stage2_f_reset_rsps$ENQ = RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    assign RTL__stage2_f_reset_rsps$DEQ = RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    assign RTL__stage2_f_reset_rsps$CLR = RTL__stage2_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__stage2_f_reset_rsps$FULL_N = RTL__stage2_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__stage2_f_reset_rsps$EMPTY_N = RTL__stage2_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    assign RTL__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__stage2_f_reset_rsps__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__stage2_f_reset_rsps__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    assign RTL__RST_N = RTL__stage3_f_reset_reqs__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    assign RTL__CLK = RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    assign RTL__stage3_f_reset_reqs$ENQ = RTL__stage3_f_reset_reqs__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    assign RTL__stage3_f_reset_reqs$FULL_N = RTL__stage3_f_reset_reqs__FULL_N;
    assign RTL__stage3_f_reset_reqs$EMPTY_N = RTL__stage3_f_reset_reqs__EMPTY_N;
    assign RTL__stage3_f_reset_reqs__RST = RTL__RST_N;
    assign RTL__stage3_f_reset_reqs__CLK = RTL__CLK;
    assign RTL__stage3_f_reset_reqs__ENQ = RTL__stage3_f_reset_reqs$ENQ;
    assign RTL__stage3_f_reset_reqs__CLR = RTL__stage3_f_reset_reqs$CLR;
    assign RTL__stage3_f_reset_rsps__DEQ = RTL__stage3_f_reset_rsps$DEQ;
    assign RTL__CLK = RTL__stage3_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__stage3_f_reset_rsps$ENQ = RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__stage3_f_reset_rsps$DEQ = RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__stage3_f_reset_rsps$CLR = RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    assign RTL__stage3_f_reset_rsps$FULL_N = RTL__stage3_f_reset_rsps__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    assign RTL__stage3_f_reset_rsps$EMPTY_N = RTL__stage3_f_reset_rsps__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    assign RTL__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__stage3_f_reset_rsps__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__stage3_f_reset_rsps__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
     
  assign  RTL__CAN_FIRE_RL_rl_show_pipe = RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL__rg_state !=4'd0&& RTL__rg_state !=4'd1&& RTL__rg_state !=4'd12; 
  assign  RTL__WILL_FIRE_RL_rl_show_pipe = RTL__CAN_FIRE_RL_rl_show_pipe ; 
  assign  RTL__CAN_FIRE_RL_rl_reset_complete = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__WILL_FIRE_RL_rl_reset_complete = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__CAN_FIRE_RL_rl_pipe = RTL__rg_state ==4'd3&&( RTL__stage3_rg_full || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0|| RTL__stage1_rg_full )&&( RTL__stage3_rg_full || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)&&( RTL__stage3_rg_full || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0||! RTL__stage1_rg_full || RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 )&&( RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0|| RTL__stage3_rg_full ); 
  assign  RTL__WILL_FIRE_RL_rl_pipe = RTL__CAN_FIRE_RL_rl_pipe ; 
  assign  RTL__CAN_FIRE_RL_rl_stage2_nonpipe = RTL__rg_state ==4'd3&&! RTL__stage3_rg_full && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3; 
  assign  RTL__WILL_FIRE_RL_rl_stage2_nonpipe = RTL__CAN_FIRE_RL_rl_stage2_nonpipe ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_trap = RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd11; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_trap = RTL__CAN_FIRE_RL_rl_stage1_trap ; 
  assign  RTL__CAN_FIRE_RL_rl_trap = RTL__rg_state ==4'd4&&(! RTL__stage1_rg_full || RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 ); 
  assign  RTL__WILL_FIRE_RL_rl_trap = RTL__CAN_FIRE_RL_rl_trap ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_CSRR_W = RTL__MUX_rg_state$write_1__SEL_9 ; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_CSRR_W = RTL__MUX_rg_state$write_1__SEL_9 ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_CSRR_W_2 = RTL__rg_state ==4'd6; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 = RTL__rg_state ==4'd6; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_CSRR_S_or_C = RTL__MUX_rg_state$write_1__SEL_10 ; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C = RTL__MUX_rg_state$write_1__SEL_10 ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_CSRR_S_or_C_2 = RTL__rg_state ==4'd7; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 = RTL__rg_state ==4'd7; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_restart_after_csrrx = RTL__rg_state ==4'd8; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx = RTL__CAN_FIRE_RL_rl_stage1_restart_after_csrrx ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_xRET = RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 &&( RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd7|| RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd8|| RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd9); 
  assign  RTL__WILL_FIRE_RL_rl_stage1_xRET = RTL__CAN_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_FENCE_I = RTL__near_mem$RDY_server_fence_i_request_put && RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd5; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_FENCE_I = RTL__CAN_FIRE_RL_rl_stage1_FENCE_I ; 
  assign  RTL__CAN_FIRE_RL_rl_finish_FENCE_I = RTL__near_mem$RDY_server_fence_i_response_get && RTL__rg_state ==4'd9; 
  assign  RTL__WILL_FIRE_RL_rl_finish_FENCE_I = RTL__CAN_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_FENCE = RTL__near_mem$RDY_server_fence_request_put && RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd4; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_FENCE = RTL__CAN_FIRE_RL_rl_stage1_FENCE ; 
  assign  RTL__CAN_FIRE_RL_rl_finish_FENCE = RTL__near_mem$RDY_server_fence_response_get && RTL__rg_state ==4'd10; 
  assign  RTL__WILL_FIRE_RL_rl_finish_FENCE = RTL__CAN_FIRE_RL_rl_finish_FENCE ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_SFENCE_VMA = RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd6; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA = RTL__CAN_FIRE_RL_rl_stage1_SFENCE_VMA ; 
  assign  RTL__CAN_FIRE_RL_rl_finish_SFENCE_VMA = RTL__rg_state ==4'd11; 
  assign  RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA = RTL__CAN_FIRE_RL_rl_finish_SFENCE_VMA ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_WFI = RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd10; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_WFI = RTL__CAN_FIRE_RL_rl_stage1_WFI ; 
  assign  RTL__CAN_FIRE_RL_rl_WFI_resume = RTL__rg_state ==4'd12&& RTL__csr_regfile$wfi_resume ; 
  assign  RTL__WILL_FIRE_RL_rl_WFI_resume = RTL__CAN_FIRE_RL_rl_WFI_resume ; 
  assign  RTL__CAN_FIRE_RL_rl_reset_from_WFI = RTL__rg_state ==4'd12&& RTL__f_reset_reqs$EMPTY_N ; 
  assign  RTL__WILL_FIRE_RL_rl_reset_from_WFI = RTL__MUX_rg_state$write_1__SEL_4 ; 
  assign  RTL__CAN_FIRE_RL_rl_trap_fetch = RTL__rg_state ==4'd5; 
  assign  RTL__WILL_FIRE_RL_rl_trap_fetch = RTL__CAN_FIRE_RL_rl_trap_fetch ; 
  assign  RTL__CAN_FIRE_RL_rl_stage1_interrupt =( RTL__csr_regfile$interrupt_pending [4]|| RTL__csr_regfile$nmi_pending )&& RTL__rg_state ==4'd3&& RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d910 && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0&&! RTL__stage3_rg_full ; 
  assign  RTL__WILL_FIRE_RL_rl_stage1_interrupt = RTL__CAN_FIRE_RL_rl_stage1_interrupt ; 
  assign  RTL__CAN_FIRE_RL_rl_reset_start = RTL__gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 && RTL__rg_state ==4'd0; 
  assign  RTL__WILL_FIRE_RL_rl_reset_start = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__CAN_FIRE_RL_stage3_rl_reset = RTL__stage3_f_reset_reqs$EMPTY_N && RTL__stage3_f_reset_rsps$FULL_N ; 
  assign  RTL__WILL_FIRE_RL_stage3_rl_reset = RTL__CAN_FIRE_RL_stage3_rl_reset ; 
  assign  RTL__CAN_FIRE_RL_stage2_rl_reset_end = RTL__stage2_f_reset_rsps$FULL_N && RTL__stage2_rg_resetting ; 
  assign  RTL__WILL_FIRE_RL_stage2_rl_reset_end = RTL__CAN_FIRE_RL_stage2_rl_reset_end ; 
  assign  RTL__CAN_FIRE_RL_stage2_rl_reset_begin = RTL__stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL__WILL_FIRE_RL_stage2_rl_reset_begin = RTL__stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL__CAN_FIRE_RL_stage1_rl_reset = RTL__stage1_f_reset_reqs$EMPTY_N && RTL__stage1_f_reset_rsps$FULL_N ; 
  assign  RTL__WILL_FIRE_RL_stage1_rl_reset = RTL__CAN_FIRE_RL_stage1_rl_reset ; 
  assign  RTL__MUX_csr_regfile$mav_csr_write_1__SEL_1 = RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 ; 
  assign  RTL__MUX_gpr_regfile$write_rd_1__SEL_3 = RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 ; 
  assign  RTL__MUX_near_mem$imem_req_1__SEL_1 = RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset ; 
  assign  RTL__MUX_near_mem$imem_req_1__SEL_2 = RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 ; 
  assign  RTL__MUX_near_mem$imem_req_1__SEL_5 = RTL__WILL_FIRE_RL_rl_WFI_resume || RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_finish_FENCE || RTL__WILL_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL__MUX_rg_next_pc$write_1__SEL_1 = RTL__WILL_FIRE_RL_rl_stage1_WFI || RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_stage1_FENCE || RTL__WILL_FIRE_RL_rl_stage1_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W ; 
  assign  RTL__MUX_rg_retiring$write_1__SEL_1 = RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2; 
  assign  RTL__MUX_rg_state$write_1__SEL_1 = RTL__gpr_regfile_RDY_server_reset_response_get__76__ETC___d688 && RTL__rg_state ==4'd1; 
  assign  RTL__MUX_rg_state$write_1__SEL_4 = RTL__CAN_FIRE_RL_rl_reset_from_WFI &&! RTL__WILL_FIRE_RL_rl_WFI_resume ; 
  assign  RTL__MUX_rg_state$write_1__SEL_6 = RTL__WILL_FIRE_RL_rl_trap_fetch || RTL__WILL_FIRE_RL_rl_WFI_resume || RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_finish_FENCE || RTL__WILL_FIRE_RL_rl_finish_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx ; 
  assign  RTL__MUX_rg_state$write_1__SEL_7 = RTL__WILL_FIRE_RL_rl_stage1_interrupt || RTL__WILL_FIRE_RL_rl_stage1_trap || RTL__WILL_FIRE_RL_rl_stage2_nonpipe ; 
  assign  RTL__MUX_rg_state$write_1__SEL_8 = RTL__WILL_FIRE_RL_rl_stage1_xRET || RTL__WILL_FIRE_RL_rl_trap ; 
  assign  RTL__MUX_rg_state$write_1__SEL_9 = RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd2; 
  assign  RTL__MUX_rg_state$write_1__SEL_10 = RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd3; 
  assign  RTL__MUX_rg_trap_info$write_1__SEL_1 = RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W ; 
  assign  RTL__MUX_rg_trap_instr$write_1__SEL_1 = RTL__WILL_FIRE_RL_rl_stage1_interrupt || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_stage1_trap ; 
  assign  RTL__MUX_rg_trap_interrupt$write_1__SEL_1 = RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_stage1_trap || RTL__WILL_FIRE_RL_rl_stage2_nonpipe ; 
  always @(     RTL__rg_trap_instr                or   RTL__csr_regfile$read_csr            or   RTL__y__h12191           or   RTL__IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868  )
         begin 
             case ( RTL__rg_trap_instr [14:12])
              3 'b010,3'b110: 
                  RTL__MUX_csr_regfile$mav_csr_write_2__VAL_2  = RTL__IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868 ;
              default : 
                  RTL__MUX_csr_regfile$mav_csr_write_2__VAL_2  = RTL__csr_regfile$read_csr [31:0]& RTL__y__h12191 ;endcase
         end
  assign  RTL__MUX_rg_state$write_1__VAL_1 = RTL__rg_run_on_reset  ? 4'd3:4'd2; 
  assign  RTL__MUX_rg_state$write_1__VAL_2 = RTL__csr_regfile$access_permitted_1  ? 4'd8:4'd4; 
  assign  RTL__MUX_rg_state$write_1__VAL_3 = RTL__csr_regfile$access_permitted_2  ? 4'd8:4'd4; 
  assign  RTL__MUX_rg_trap_info$write_1__VAL_1 ={ RTL__near_mem$imem_pc ,4'd2, RTL__value__h6967 }; 
  assign  RTL__MUX_rg_trap_info$write_1__VAL_2 ={ RTL__stage2_rg_stage2 [166:135], RTL__near_mem$dmem_exc_code , RTL__stage2_rg_stage2 [95:64]}; 
  assign  RTL__MUX_rg_trap_info$write_1__VAL_3 ={ RTL__near_mem$imem_pc , RTL__IF_near_mem_imem_exc__78_THEN_near_mem_imem_ex_ETC___d799 }; 
  assign  RTL__MUX_rg_trap_info$write_1__VAL_4 ={ RTL__near_mem$imem_pc , RTL__x_exc_code__h15410 ,32'd0}; 
  assign  RTL__MUX_s1_to_s2$write_1__VAL_1 = RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ; 
  assign  RTL__MUX_stage1_rg_full$write_1__VAL_10 = RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d776 ||( RTL__csr_regfile_interrupt_pending_rg_cur_priv_9_07_ETC___d779 || RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 )&& RTL__stage1_rg_full ; 
  assign  RTL__MUX_stage2_rg_full$write_1__VAL_3 = RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d769 || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd2&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0; 
  assign  RTL__cfg_logdelay$D_IN = RTL__set_verbosity_logdelay ; 
  assign  RTL__cfg_logdelay$EN = RTL__EN_set_verbosity ; 
  assign  RTL__cfg_verbosity$D_IN = RTL__set_verbosity_verbosity ; 
  assign  RTL__cfg_verbosity$EN = RTL__EN_set_verbosity ; 
  assign  RTL__rg_csr_pc$D_IN = RTL__near_mem$imem_pc ; 
  assign  RTL__rg_csr_pc$EN = RTL__MUX_rg_trap_info$write_1__SEL_1 ; 
  assign  RTL__rg_csr_val1$D_IN = RTL__x_out_data_to_stage2_val1__h5224 ; 
  assign  RTL__rg_csr_val1$EN = RTL__MUX_rg_trap_info$write_1__SEL_1 ; 
  always @(      RTL__WILL_FIRE_RL_rl_trap                  or   RTL__csr_regfile$csr_trap_actions             or   RTL__WILL_FIRE_RL_rl_stage1_xRET            or   RTL__csr_regfile$csr_ret_actions           or   RTL__WILL_FIRE_RL_rl_reset_start  )
         begin 
             case (1'b1) 
              RTL__WILL_FIRE_RL_rl_trap  : 
                  RTL__rg_cur_priv$D_IN  = RTL__csr_regfile$csr_trap_actions [1:0]; 
              RTL__WILL_FIRE_RL_rl_stage1_xRET  : 
                  RTL__rg_cur_priv$D_IN  = RTL__csr_regfile$csr_ret_actions [33:32]; 
              RTL__WILL_FIRE_RL_rl_reset_start  : 
                  RTL__rg_cur_priv$D_IN  =2'b11;
              default : 
                  RTL__rg_cur_priv$D_IN  =2'b10;endcase
         end
  assign  RTL__rg_cur_priv$EN = RTL__WILL_FIRE_RL_rl_trap || RTL__WILL_FIRE_RL_rl_stage1_xRET || RTL__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__rg_mstatus_MXR$D_IN = RTL__csr_regfile$read_mstatus [19]; 
  assign  RTL__rg_mstatus_MXR$EN = RTL__MUX_rg_state$write_1__SEL_8 ; 
  always @(       RTL__MUX_rg_next_pc$write_1__SEL_1                    or   RTL__x_out_next_pc__h5189              or   RTL__WILL_FIRE_RL_rl_trap             or   RTL__csr_regfile$csr_trap_actions            or   RTL__WILL_FIRE_RL_rl_stage1_xRET           or   RTL__csr_regfile$csr_ret_actions  )
         begin 
             case (1'b1) 
              RTL__MUX_rg_next_pc$write_1__SEL_1  : 
                  RTL__rg_next_pc$D_IN  = RTL__x_out_next_pc__h5189 ; 
              RTL__WILL_FIRE_RL_rl_trap  : 
                  RTL__rg_next_pc$D_IN  = RTL__csr_regfile$csr_trap_actions [97:66]; 
              RTL__WILL_FIRE_RL_rl_stage1_xRET  : 
                  RTL__rg_next_pc$D_IN  = RTL__csr_regfile$csr_ret_actions [65:34];
              default : 
                  RTL__rg_next_pc$D_IN  =32'hAAAAAAAA;endcase
         end
  assign  RTL__rg_next_pc$EN = RTL__WILL_FIRE_RL_rl_stage1_WFI || RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_stage1_FENCE || RTL__WILL_FIRE_RL_rl_stage1_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_trap || RTL__WILL_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL__rg_retiring$D_IN =1'd1; 
  assign  RTL__rg_retiring$EN = RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 || RTL__WILL_FIRE_RL_rl_stage1_WFI || RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_stage1_FENCE || RTL__WILL_FIRE_RL_rl_stage1_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_xRET || RTL__WILL_FIRE_RL_rl_trap || RTL__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__rg_run_on_reset$D_IN = RTL__f_reset_reqs$D_OUT ; 
  assign  RTL__rg_run_on_reset$EN = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__rg_sstatus_SUM$D_IN =1'd0; 
  assign  RTL__rg_sstatus_SUM$EN = RTL__MUX_rg_state$write_1__SEL_8 ; 
  assign  RTL__rg_start_CPI_cycles$D_IN = RTL__csr_regfile$read_csr_mcycle ; 
  assign  RTL__rg_start_CPI_cycles$EN = RTL__MUX_near_mem$imem_req_1__SEL_1 ; 
  assign  RTL__rg_start_CPI_instrs$D_IN = RTL__csr_regfile$read_csr_minstret ; 
  assign  RTL__rg_start_CPI_instrs$EN = RTL__MUX_near_mem$imem_req_1__SEL_1 ; 
  always @(                  RTL__WILL_FIRE_RL_rl_reset_complete                                          or   RTL__MUX_rg_state$write_1__VAL_1                         or   RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2                        or   RTL__MUX_rg_state$write_1__VAL_2                       or   RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2                      or   RTL__MUX_rg_state$write_1__VAL_3                     or   RTL__WILL_FIRE_RL_rl_reset_from_WFI                    or   RTL__WILL_FIRE_RL_rl_reset_start                   or   RTL__MUX_rg_state$write_1__SEL_6                  or   RTL__MUX_rg_state$write_1__SEL_7                 or   RTL__MUX_rg_state$write_1__SEL_8                or   RTL__WILL_FIRE_RL_rl_stage1_CSRR_W               or   RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C              or   RTL__WILL_FIRE_RL_rl_stage1_FENCE_I             or   RTL__WILL_FIRE_RL_rl_stage1_FENCE            or   RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA           or   RTL__WILL_FIRE_RL_rl_stage1_WFI  )
         begin 
             case (1'b1) 
              RTL__WILL_FIRE_RL_rl_reset_complete  : 
                  RTL__rg_state$D_IN  = RTL__MUX_rg_state$write_1__VAL_1 ; 
              RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2  : 
                  RTL__rg_state$D_IN  = RTL__MUX_rg_state$write_1__VAL_2 ; 
              RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2  : 
                  RTL__rg_state$D_IN  = RTL__MUX_rg_state$write_1__VAL_3 ; 
              RTL__WILL_FIRE_RL_rl_reset_from_WFI  : 
                  RTL__rg_state$D_IN  =4'd0; 
              RTL__WILL_FIRE_RL_rl_reset_start  : 
                  RTL__rg_state$D_IN  =4'd1; 
              RTL__MUX_rg_state$write_1__SEL_6  : 
                  RTL__rg_state$D_IN  =4'd3; 
              RTL__MUX_rg_state$write_1__SEL_7  : 
                  RTL__rg_state$D_IN  =4'd4; 
              RTL__MUX_rg_state$write_1__SEL_8  : 
                  RTL__rg_state$D_IN  =4'd5; 
              RTL__WILL_FIRE_RL_rl_stage1_CSRR_W  : 
                  RTL__rg_state$D_IN  =4'd6; 
              RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C  : 
                  RTL__rg_state$D_IN  =4'd7; 
              RTL__WILL_FIRE_RL_rl_stage1_FENCE_I  : 
                  RTL__rg_state$D_IN  =4'd9; 
              RTL__WILL_FIRE_RL_rl_stage1_FENCE  : 
                  RTL__rg_state$D_IN  =4'd10; 
              RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA  : 
                  RTL__rg_state$D_IN  =4'd11; 
              RTL__WILL_FIRE_RL_rl_stage1_WFI  : 
                  RTL__rg_state$D_IN  =4'd12;
              default : 
                  RTL__rg_state$D_IN  =4'b1010;endcase
         end
  assign  RTL__rg_state$EN = RTL__WILL_FIRE_RL_rl_reset_complete || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 || RTL__WILL_FIRE_RL_rl_reset_from_WFI || RTL__WILL_FIRE_RL_rl_reset_start || RTL__WILL_FIRE_RL_rl_trap_fetch || RTL__WILL_FIRE_RL_rl_WFI_resume || RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_finish_FENCE || RTL__WILL_FIRE_RL_rl_finish_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx || RTL__WILL_FIRE_RL_rl_stage1_interrupt || RTL__WILL_FIRE_RL_rl_stage1_trap || RTL__WILL_FIRE_RL_rl_stage2_nonpipe || RTL__WILL_FIRE_RL_rl_stage1_xRET || RTL__WILL_FIRE_RL_rl_trap || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_FENCE || RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_stage1_WFI ; 
  always @(         RTL__MUX_rg_trap_info$write_1__SEL_1                        or   RTL__MUX_rg_trap_info$write_1__VAL_1                or   RTL__WILL_FIRE_RL_rl_stage2_nonpipe               or   RTL__MUX_rg_trap_info$write_1__VAL_2              or   RTL__WILL_FIRE_RL_rl_stage1_trap             or   RTL__MUX_rg_trap_info$write_1__VAL_3            or   RTL__WILL_FIRE_RL_rl_stage1_interrupt           or   RTL__MUX_rg_trap_info$write_1__VAL_4  )
         begin 
             case (1'b1) 
              RTL__MUX_rg_trap_info$write_1__SEL_1  : 
                  RTL__rg_trap_info$D_IN  = RTL__MUX_rg_trap_info$write_1__VAL_1 ; 
              RTL__WILL_FIRE_RL_rl_stage2_nonpipe  : 
                  RTL__rg_trap_info$D_IN  = RTL__MUX_rg_trap_info$write_1__VAL_2 ; 
              RTL__WILL_FIRE_RL_rl_stage1_trap  : 
                  RTL__rg_trap_info$D_IN  = RTL__MUX_rg_trap_info$write_1__VAL_3 ; 
              RTL__WILL_FIRE_RL_rl_stage1_interrupt  : 
                  RTL__rg_trap_info$D_IN  = RTL__MUX_rg_trap_info$write_1__VAL_4 ;
              default : 
                  RTL__rg_trap_info$D_IN  =68'hAAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL__rg_trap_info$EN = RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_stage2_nonpipe || RTL__WILL_FIRE_RL_rl_stage1_trap || RTL__WILL_FIRE_RL_rl_stage1_interrupt ; 
  assign  RTL__rg_trap_instr$D_IN = RTL__MUX_rg_trap_instr$write_1__SEL_1  ?  RTL__near_mem$imem_instr : RTL__stage2_rg_stage2 [134:103]; 
  assign  RTL__rg_trap_instr$EN = RTL__WILL_FIRE_RL_rl_stage1_interrupt || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_stage1_trap || RTL__WILL_FIRE_RL_rl_stage2_nonpipe ; 
  assign  RTL__rg_trap_interrupt$D_IN =! RTL__MUX_rg_trap_interrupt$write_1__SEL_1 ; 
  assign  RTL__rg_trap_interrupt$EN = RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL__WILL_FIRE_RL_rl_stage1_CSRR_W || RTL__WILL_FIRE_RL_rl_stage1_trap || RTL__WILL_FIRE_RL_rl_stage2_nonpipe || RTL__WILL_FIRE_RL_rl_stage1_interrupt ; 
  assign  RTL__s1_to_s2$D_IN = RTL__WILL_FIRE_RL_rl_pipe && RTL__MUX_s1_to_s2$write_1__VAL_1 ; 
  assign  RTL__s1_to_s2$EN = RTL__WILL_FIRE_RL_rl_pipe || RTL__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__s2_to_s3$D_IN = RTL__MUX_rg_retiring$write_1__SEL_1 ; 
  assign  RTL__s2_to_s3$EN = RTL__WILL_FIRE_RL_rl_pipe || RTL__WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL__s3_deq$D_IN = RTL__WILL_FIRE_RL_rl_pipe && RTL__stage3_rg_full ; 
  assign  RTL__s3_deq$EN = RTL__WILL_FIRE_RL_rl_pipe || RTL__WILL_FIRE_RL_rl_reset_start ; 
  always @(             RTL__WILL_FIRE_RL_stage1_rl_reset                                or   RTL__WILL_FIRE_RL_rl_trap_fetch                    or   RTL__WILL_FIRE_RL_rl_WFI_resume                   or   RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA                  or   RTL__WILL_FIRE_RL_rl_finish_FENCE                 or   RTL__WILL_FIRE_RL_rl_finish_FENCE_I                or   RTL__WILL_FIRE_RL_rl_stage1_xRET               or   RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx              or   RTL__WILL_FIRE_RL_rl_trap             or   RTL__WILL_FIRE_RL_rl_pipe            or   RTL__MUX_stage1_rg_full$write_1__VAL_10           or   RTL__MUX_near_mem$imem_req_1__SEL_1  )
         case (1'b1) 
          RTL__WILL_FIRE_RL_stage1_rl_reset  : 
              RTL__stage1_rg_full$D_IN  =1'd0; 
          RTL__WILL_FIRE_RL_rl_trap_fetch  || RTL__WILL_FIRE_RL_rl_WFI_resume || RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_finish_FENCE || RTL__WILL_FIRE_RL_rl_finish_FENCE_I : 
              RTL__stage1_rg_full$D_IN  =1'd1; 
          RTL__WILL_FIRE_RL_rl_stage1_xRET  : 
              RTL__stage1_rg_full$D_IN  =1'd0; 
          RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx  : 
              RTL__stage1_rg_full$D_IN  =1'd1; 
          RTL__WILL_FIRE_RL_rl_trap  : 
              RTL__stage1_rg_full$D_IN  =1'd0; 
          RTL__WILL_FIRE_RL_rl_pipe  : 
              RTL__stage1_rg_full$D_IN  = RTL__MUX_stage1_rg_full$write_1__VAL_10 ; 
          RTL__MUX_near_mem$imem_req_1__SEL_1  : 
              RTL__stage1_rg_full$D_IN  =1'd1;
          default : 
              RTL__stage1_rg_full$D_IN  =1'b0;endcase
  assign  RTL__stage1_rg_full$EN = RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset || RTL__WILL_FIRE_RL_rl_pipe || RTL__WILL_FIRE_RL_rl_stage1_xRET || RTL__WILL_FIRE_RL_rl_trap || RTL__WILL_FIRE_RL_stage1_rl_reset || RTL__WILL_FIRE_RL_rl_trap_fetch || RTL__WILL_FIRE_RL_rl_WFI_resume || RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_finish_FENCE || RTL__WILL_FIRE_RL_rl_finish_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx ; 
  always @(      RTL__stage2_f_reset_reqs$EMPTY_N                  or   RTL__WILL_FIRE_RL_rl_trap             or   RTL__WILL_FIRE_RL_rl_pipe            or   RTL__MUX_stage2_rg_full$write_1__VAL_3           or   RTL__MUX_near_mem$imem_req_1__SEL_1  )
         case (1'b1) 
          RTL__stage2_f_reset_reqs$EMPTY_N  || RTL__WILL_FIRE_RL_rl_trap : 
              RTL__stage2_rg_full$D_IN  =1'd0; 
          RTL__WILL_FIRE_RL_rl_pipe  : 
              RTL__stage2_rg_full$D_IN  = RTL__MUX_stage2_rg_full$write_1__VAL_3 ; 
          RTL__MUX_near_mem$imem_req_1__SEL_1  : 
              RTL__stage2_rg_full$D_IN  =1'd0;
          default : 
              RTL__stage2_rg_full$D_IN  =1'b0;endcase
  assign  RTL__stage2_rg_full$EN = RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset || RTL__WILL_FIRE_RL_rl_pipe || RTL__WILL_FIRE_RL_rl_trap || RTL__stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL__stage2_rg_resetting$D_IN = RTL__stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL__stage2_rg_resetting$EN = RTL__WILL_FIRE_RL_stage2_rl_reset_end || RTL__stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL__stage2_rg_stage2$D_IN ={ RTL__rg_cur_priv , RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 , RTL__x_out_data_to_stage2_rd__h5222 , RTL__x_out_data_to_stage2_addr__h5223 , RTL__x_out_data_to_stage2_val1__h5224 , RTL__x_out_data_to_stage2_val2__h5225 }; 
  assign  RTL__stage2_rg_stage2$EN = RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 ; 
  always @(     RTL__WILL_FIRE_RL_stage3_rl_reset                or   RTL__WILL_FIRE_RL_rl_pipe            or   RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86           or   RTL__MUX_near_mem$imem_req_1__SEL_1  )
         case (1'b1) 
          RTL__WILL_FIRE_RL_stage3_rl_reset  : 
              RTL__stage3_rg_full$D_IN  =1'd0; 
          RTL__WILL_FIRE_RL_rl_pipe  : 
              RTL__stage3_rg_full$D_IN  = RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2; 
          RTL__MUX_near_mem$imem_req_1__SEL_1  : 
              RTL__stage3_rg_full$D_IN  =1'd0;
          default : 
              RTL__stage3_rg_full$D_IN  =1'b0;endcase
  assign  RTL__stage3_rg_full$EN = RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset || RTL__WILL_FIRE_RL_rl_pipe || RTL__WILL_FIRE_RL_stage3_rl_reset ; 
  assign  RTL__stage3_rg_stage3$D_IN ={ RTL__stage2_rg_stage2 [166:103], RTL__stage2_rg_stage2 [168:167], RTL__stage2_rg_stage2 [102:101]==2'd0|| RTL__near_mem$dmem_valid &&! RTL__near_mem$dmem_exc , RTL__x_out_data_to_stage3_rd__h4667 , RTL__x_out_data_to_stage3_rd_val__h4668 }; 
  assign  RTL__stage3_rg_stage3$EN = RTL__MUX_rg_retiring$write_1__SEL_1 ; 
  assign  RTL__csr_regfile$access_permitted_1_csr_addr = RTL__rg_trap_instr [31:20]; 
  assign  RTL__csr_regfile$access_permitted_1_priv = RTL__rg_cur_priv ; 
  assign  RTL__csr_regfile$access_permitted_1_read_not_write =1'd0; 
  assign  RTL__csr_regfile$access_permitted_2_csr_addr = RTL__rg_trap_instr [31:20]; 
  assign  RTL__csr_regfile$access_permitted_2_priv = RTL__rg_cur_priv ; 
  assign  RTL__csr_regfile$access_permitted_2_read_not_write = RTL__rs1_val__h11920 ==32'd0; 
  assign  RTL__csr_regfile$csr_counter_read_fault_csr_addr =12'h0; 
  assign  RTL__csr_regfile$csr_counter_read_fault_priv =2'h0; 
  always @(  RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415  )
         begin 
             case ( RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 )
              4 'd7: 
                  RTL__csr_regfile$csr_ret_actions_from_priv  =2'b11;
              4 'd8: 
                  RTL__csr_regfile$csr_ret_actions_from_priv  =2'b01;
              default : 
                  RTL__csr_regfile$csr_ret_actions_from_priv  =2'b0;endcase
         end
  assign  RTL__csr_regfile$csr_trap_actions_exc_code = RTL__rg_trap_info [35:32]; 
  assign  RTL__csr_regfile$csr_trap_actions_from_priv = RTL__rg_cur_priv ; 
  assign  RTL__csr_regfile$csr_trap_actions_interrupt = RTL__rg_trap_interrupt &&! RTL__csr_regfile$nmi_pending ; 
  assign  RTL__csr_regfile$csr_trap_actions_nmi = RTL__rg_trap_interrupt && RTL__csr_regfile$nmi_pending ; 
  assign  RTL__csr_regfile$csr_trap_actions_pc = RTL__rg_trap_info [67:36]; 
  assign  RTL__csr_regfile$csr_trap_actions_xtval = RTL__rg_trap_info [31:0]; 
  assign  RTL__csr_regfile$interrupt_pending_cur_priv = RTL__rg_cur_priv ; 
  assign  RTL__csr_regfile$m_external_interrupt_req_set_not_clear = RTL__m_external_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile$mav_csr_write_csr_addr = RTL__rg_trap_instr [31:20]; 
  assign  RTL__csr_regfile$mav_csr_write_word = RTL__MUX_csr_regfile$mav_csr_write_1__SEL_1  ?  RTL__rs1_val__h11213 : RTL__MUX_csr_regfile$mav_csr_write_2__VAL_2 ; 
  assign  RTL__csr_regfile$mav_read_csr_csr_addr =12'h0; 
  assign  RTL__csr_regfile$nmi_req_set_not_clear = RTL__nmi_req_set_not_clear ; 
  assign  RTL__csr_regfile$read_csr_csr_addr = RTL__rg_trap_instr [31:20]; 
  assign  RTL__csr_regfile$read_csr_port2_csr_addr =12'h0; 
  assign  RTL__csr_regfile$s_external_interrupt_req_set_not_clear = RTL__s_external_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile$software_interrupt_req_set_not_clear = RTL__software_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile$timer_interrupt_req_set_not_clear = RTL__timer_interrupt_req_set_not_clear ; 
  assign  RTL__csr_regfile$EN_server_reset_request_put = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__csr_regfile$EN_server_reset_response_get = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__csr_regfile$EN_mav_read_csr =1'b0; 
  assign  RTL__csr_regfile$EN_mav_csr_write = RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 && RTL__rg_trap_instr [19:15]!=5'd0; 
  assign  RTL__csr_regfile$EN_csr_trap_actions = RTL__CAN_FIRE_RL_rl_trap ; 
  assign  RTL__csr_regfile$EN_csr_ret_actions = RTL__CAN_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL__csr_regfile$EN_csr_minstret_incr = RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 || RTL__WILL_FIRE_RL_rl_stage1_WFI || RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_stage1_FENCE || RTL__WILL_FIRE_RL_rl_stage1_FENCE_I || RTL__WILL_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL__csr_regfile$EN_debug =1'b0; 
  assign  RTL__f_reset_reqs$D_IN = RTL__hart0_server_reset_request_put ; 
  assign  RTL__f_reset_reqs$ENQ = RTL__EN_hart0_server_reset_request_put ; 
  assign  RTL__f_reset_reqs$DEQ = RTL__gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 && RTL__rg_state ==4'd0; 
  assign  RTL__f_reset_reqs$CLR =1'b0; 
  assign  RTL__f_reset_rsps$D_IN = RTL__rg_run_on_reset ; 
  assign  RTL__f_reset_rsps$ENQ = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__f_reset_rsps$DEQ = RTL__EN_hart0_server_reset_response_get ; 
  assign  RTL__f_reset_rsps$CLR =1'b0; 
  assign  RTL__gpr_regfile$read_rs1_port2_rs1 =5'h0; 
  assign  RTL__gpr_regfile$read_rs1_rs1 = RTL__near_mem$imem_instr [19:15]; 
  assign  RTL__gpr_regfile$read_rs2_rs2 = RTL__near_mem$imem_instr [24:20]; 
  assign  RTL__gpr_regfile$write_rd_rd =( RTL__MUX_csr_regfile$mav_csr_write_1__SEL_1 || RTL__MUX_gpr_regfile$write_rd_1__SEL_3 ) ?  RTL__rg_trap_instr [11:7]: RTL__stage3_rg_stage3 [36:32]; 
  assign  RTL__gpr_regfile$write_rd_rd_val =( RTL__MUX_csr_regfile$mav_csr_write_1__SEL_1 || RTL__MUX_gpr_regfile$write_rd_1__SEL_3 ) ?  RTL__csr_regfile$read_csr [31:0]: RTL__stage3_rg_stage3 [31:0]; 
  assign  RTL__gpr_regfile$EN_server_reset_request_put = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__gpr_regfile$EN_server_reset_response_get = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__gpr_regfile$EN_write_rd = RTL__WILL_FIRE_RL_rl_pipe && RTL__stage3_rg_full && RTL__stage3_rg_stage3 [37]|| RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 || RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 ; 
  assign  RTL__near_mem$dmem_master_arready = RTL__dmem_master_arready ; 
  assign  RTL__near_mem$dmem_master_awready = RTL__dmem_master_awready ; 
  assign  RTL__near_mem$dmem_master_bid = RTL__dmem_master_bid ; 
  assign  RTL__near_mem$dmem_master_bresp = RTL__dmem_master_bresp ; 
  assign  RTL__near_mem$dmem_master_bvalid = RTL__dmem_master_bvalid ; 
  assign  RTL__near_mem$dmem_master_rdata = RTL__dmem_master_rdata ; 
  assign  RTL__near_mem$dmem_master_rid = RTL__dmem_master_rid ; 
  assign  RTL__near_mem$dmem_master_rlast = RTL__dmem_master_rlast ; 
  assign  RTL__near_mem$dmem_master_rresp = RTL__dmem_master_rresp ; 
  assign  RTL__near_mem$dmem_master_rvalid = RTL__dmem_master_rvalid ; 
  assign  RTL__near_mem$dmem_master_wready = RTL__dmem_master_wready ; 
  assign  RTL__near_mem$dmem_req_addr = RTL__x_out_data_to_stage2_addr__h5223 ; 
  assign  RTL__near_mem$dmem_req_f3 = RTL__near_mem$imem_instr [14:12]; 
  assign  RTL__near_mem$dmem_req_mstatus_MXR = RTL__csr_regfile$read_mstatus [19]; 
  assign  RTL__near_mem$dmem_req_op = RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd1; 
  assign  RTL__near_mem$dmem_req_priv = RTL__csr_regfile$read_mstatus [17] ?  RTL__csr_regfile$read_mstatus [12:11]: RTL__rg_cur_priv ; 
  assign  RTL__near_mem$dmem_req_satp = RTL__csr_regfile$read_satp ; 
  assign  RTL__near_mem$dmem_req_sstatus_SUM =1'd0; 
  assign  RTL__near_mem$dmem_req_store_value ={32'd0, RTL__x_out_data_to_stage2_val2__h5225 }; 
  assign  RTL__near_mem$imem_master_arready = RTL__imem_master_arready ; 
  assign  RTL__near_mem$imem_master_awready = RTL__imem_master_awready ; 
  assign  RTL__near_mem$imem_master_bid = RTL__imem_master_bid ; 
  assign  RTL__near_mem$imem_master_bresp = RTL__imem_master_bresp ; 
  assign  RTL__near_mem$imem_master_bvalid = RTL__imem_master_bvalid ; 
  assign  RTL__near_mem$imem_master_rdata = RTL__imem_master_rdata ; 
  assign  RTL__near_mem$imem_master_rid = RTL__imem_master_rid ; 
  assign  RTL__near_mem$imem_master_rlast = RTL__imem_master_rlast ; 
  assign  RTL__near_mem$imem_master_rresp = RTL__imem_master_rresp ; 
  assign  RTL__near_mem$imem_master_rvalid = RTL__imem_master_rvalid ; 
  assign  RTL__near_mem$imem_master_wready = RTL__imem_master_wready ; 
  always @(         RTL__MUX_near_mem$imem_req_1__SEL_1                        or   RTL__soc_map$m_pc_reset_value                or   RTL__WILL_FIRE_RL_rl_trap_fetch               or   RTL__MUX_near_mem$imem_req_1__SEL_5              or   RTL__rg_next_pc             or   RTL__MUX_near_mem$imem_req_1__SEL_2            or   RTL__x_out_next_pc__h5189           or   RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx  )
         begin 
             case (1'b1) 
              RTL__MUX_near_mem$imem_req_1__SEL_1  : 
                  RTL__near_mem$imem_req_addr  = RTL__soc_map$m_pc_reset_value [31:0]; 
              RTL__WILL_FIRE_RL_rl_trap_fetch  || RTL__MUX_near_mem$imem_req_1__SEL_5 : 
                  RTL__near_mem$imem_req_addr  = RTL__rg_next_pc ; 
              RTL__MUX_near_mem$imem_req_1__SEL_2  : 
                  RTL__near_mem$imem_req_addr  = RTL__x_out_next_pc__h5189 ; 
              RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx  : 
                  RTL__near_mem$imem_req_addr  = RTL__x_out_next_pc__h5189 ;
              default : 
                  RTL__near_mem$imem_req_addr  =32'hAAAAAAAA;endcase
         end
  assign  RTL__near_mem$imem_req_f3 =3'b010; 
  assign  RTL__near_mem$imem_req_mstatus_MXR =( RTL__MUX_near_mem$imem_req_1__SEL_1 || RTL__MUX_near_mem$imem_req_1__SEL_2 || RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx || RTL__MUX_near_mem$imem_req_1__SEL_5 ) ?  RTL__csr_regfile$read_mstatus [19]: RTL__rg_mstatus_MXR ; 
  assign  RTL__near_mem$imem_req_priv = RTL__rg_cur_priv ; 
  assign  RTL__near_mem$imem_req_satp = RTL__csr_regfile$read_satp ; 
  assign  RTL__near_mem$imem_req_sstatus_SUM = RTL__WILL_FIRE_RL_rl_trap_fetch && RTL__rg_sstatus_SUM ; 
  assign  RTL__near_mem$server_fence_request_put =8'b10101010; 
  assign  RTL__near_mem$EN_server_reset_request_put = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__near_mem$EN_server_reset_response_get = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__near_mem$EN_imem_req = RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset || RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 || RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx || RTL__WILL_FIRE_RL_rl_trap_fetch || RTL__WILL_FIRE_RL_rl_WFI_resume || RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL__WILL_FIRE_RL_rl_finish_FENCE || RTL__WILL_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL__near_mem$EN_dmem_req = RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 &&( RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd1|| RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd2); 
  assign  RTL__near_mem$EN_server_fence_i_request_put = RTL__CAN_FIRE_RL_rl_stage1_FENCE_I ; 
  assign  RTL__near_mem$EN_server_fence_i_response_get = RTL__CAN_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL__near_mem$EN_server_fence_request_put = RTL__CAN_FIRE_RL_rl_stage1_FENCE ; 
  assign  RTL__near_mem$EN_server_fence_response_get = RTL__CAN_FIRE_RL_rl_finish_FENCE ; 
  assign  RTL__near_mem$EN_sfence_vma = RTL__CAN_FIRE_RL_rl_stage1_SFENCE_VMA ; 
  assign  RTL__soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL__soc_map$m_is_mem_addr_addr =64'h0; 
  assign  RTL__soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL__stage1_f_reset_reqs$ENQ = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__stage1_f_reset_reqs$DEQ = RTL__CAN_FIRE_RL_stage1_rl_reset ; 
  assign  RTL__stage1_f_reset_reqs$CLR =1'b0; 
  assign  RTL__stage1_f_reset_rsps$ENQ = RTL__CAN_FIRE_RL_stage1_rl_reset ; 
  assign  RTL__stage1_f_reset_rsps$DEQ = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__stage1_f_reset_rsps$CLR =1'b0; 
  assign  RTL__stage2_f_reset_reqs$ENQ = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__stage2_f_reset_reqs$DEQ = RTL__stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL__stage2_f_reset_reqs$CLR =1'b0; 
  assign  RTL__stage2_f_reset_rsps$ENQ = RTL__CAN_FIRE_RL_stage2_rl_reset_end ; 
  assign  RTL__stage2_f_reset_rsps$DEQ = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__stage2_f_reset_rsps$CLR =1'b0; 
  assign  RTL__stage3_f_reset_reqs$ENQ = RTL__CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL__stage3_f_reset_reqs$DEQ = RTL__CAN_FIRE_RL_stage3_rl_reset ; 
  assign  RTL__stage3_f_reset_reqs$CLR =1'b0; 
  assign  RTL__stage3_f_reset_rsps$ENQ = RTL__CAN_FIRE_RL_stage3_rl_reset ; 
  assign  RTL__stage3_f_reset_rsps$DEQ = RTL__MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL__stage3_f_reset_rsps$CLR =1'b0; 
  assign  RTL__IF_IF_near_mem_imem_instr__59_BITS_6_TO_0_79_E_ETC___d655 =(( RTL__near_mem$imem_instr [6:0]==7'b1100011) ?  RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616 : RTL__near_mem$imem_instr [6:0]==7'b1101111|| RTL__near_mem$imem_instr [6:0]==7'b1100111) ?  RTL__data_to_stage2_addr__h5215 :(( RTL__near_mem$imem_instr [6:0]==7'b1110011&& RTL__near_mem$imem_instr [14:12]==3'b0&& RTL__near_mem$imem_instr [11:7]==5'd0&& RTL__near_mem$imem_instr [19:15]==5'd0&& RTL__near_mem$imem_instr [31:20]==12'b000000000001) ?  RTL__near_mem$imem_pc :32'd0); 
  assign  RTL__IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362 = RTL__NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252  ? 4'd11:4'd0; 
  assign  RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 = RTL__near_mem$imem_exc  ? 4'd11: RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413 ; 
  assign  RTL__IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868 = RTL__csr_regfile$read_csr [31:0]| RTL__rs1_val__h11920 ; 
  assign  RTL__IF_near_mem_imem_exc__78_THEN_near_mem_imem_ex_ETC___d799 = RTL__near_mem$imem_exc  ? { RTL__near_mem$imem_exc_code , RTL__near_mem$imem_tval }:{ RTL__alu_outputs_exc_code__h5862 , RTL__trap_info_tval__h6925 }; 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285 = RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 && RTL__alu_outputs___1_val2__h5367 [1]|| RTL__near_mem$imem_instr [14:12]!=3'b0&& RTL__near_mem$imem_instr [14:12]!=3'b001&& RTL__near_mem$imem_instr [14:12]!=3'b100&& RTL__near_mem$imem_instr [14:12]!=3'b101&& RTL__near_mem$imem_instr [14:12]!=3'b110&& RTL__near_mem$imem_instr [14:12]!=3'b111; 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 = RTL__rs1_val_bypassed__h3337 == RTL__rs2_val__h5339 ; 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 =( RTL__rs1_val_bypassed__h3337 ^32'h80000000)<( RTL__rs2_val__h5339 ^32'h80000000); 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 = RTL__rs1_val_bypassed__h3337 < RTL__rs2_val__h5339 ; 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 =( RTL__near_mem$imem_instr [6:0]==7'b1100011) ?  RTL__near_mem$imem_instr [14:12]!=3'b0&& RTL__near_mem$imem_instr [14:12]!=3'b001&& RTL__near_mem$imem_instr [14:12]!=3'b100&& RTL__near_mem$imem_instr [14:12]!=3'b101&& RTL__near_mem$imem_instr [14:12]!=3'b110&& RTL__near_mem$imem_instr [14:12]!=3'b111|| RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 :((( RTL__near_mem$imem_instr [6:0]==7'b0010011|| RTL__near_mem$imem_instr [6:0]==7'b0110011)&&( RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b101)) ?  RTL__near_mem$imem_instr [25]: RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8 ); 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 =( RTL__near_mem$imem_instr [6:0]==7'b1100011) ? ( RTL__near_mem$imem_instr [14:12]==3'b0|| RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b100|| RTL__near_mem$imem_instr [14:12]==3'b101|| RTL__near_mem$imem_instr [14:12]==3'b110|| RTL__near_mem$imem_instr [14:12]==3'b111)&& RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 :((( RTL__near_mem$imem_instr [6:0]==7'b0010011|| RTL__near_mem$imem_instr [6:0]==7'b0110011)&&( RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b101)) ? ! RTL__near_mem$imem_instr [25]: RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9 ); 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571 =(( RTL__near_mem$imem_instr [6:0]==7'b0010011|| RTL__near_mem$imem_instr [6:0]==7'b0110011)&&( RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b101)) ?  RTL__alu_outputs___1_val1__h5480 : RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570 ; 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d649 =( RTL__near_mem$imem_instr [6:0]==7'b1100011) ?  RTL__near_mem$imem_instr [14:12]!=3'b0&& RTL__near_mem$imem_instr [14:12]!=3'b001&& RTL__near_mem$imem_instr [14:12]!=3'b100&& RTL__near_mem$imem_instr [14:12]!=3'b101&& RTL__near_mem$imem_instr [14:12]!=3'b110&& RTL__near_mem$imem_instr [14:12]!=3'b111|| RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 ||! RTL__alu_outputs___1_val2__h5367 [1]: RTL__near_mem$imem_instr [6:0]!=7'b1101111&& RTL__near_mem$imem_instr [6:0]!=7'b1100111&&( RTL__near_mem$imem_instr [6:0]!=7'b1110011|| RTL__near_mem$imem_instr [14:12]!=3'b0|| RTL__near_mem$imem_instr [11:7]!=5'd0|| RTL__near_mem$imem_instr [19:15]!=5'd0|| RTL__near_mem$imem_instr [31:20]!=12'b0&& RTL__near_mem$imem_instr [31:20]!=12'b000000000001); 
  assign  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d910 = RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 || RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL__IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394 =(( RTL__rg_cur_priv ==2'b11|| RTL__rg_cur_priv ==2'b01&&! RTL__csr_regfile$read_mstatus [22])&& RTL__near_mem$imem_instr [31:20]==12'b000100000010) ? 4'd8:( RTL__rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_EQ_0_ETC___d392  ? 4'd10:4'd11); 
  assign  RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 = RTL__stage2_rg_full  ?  RTL__CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5 :2'd0; 
  assign  RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 = RTL__stage2_rg_stage2 [100:96]== RTL__near_mem$imem_instr [19:15]; 
  assign  RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 = RTL__stage2_rg_stage2 [100:96]== RTL__near_mem$imem_instr [24:20]; 
  assign  RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 = RTL__stage2_rg_full  ?  RTL__IF_stage2_rg_stage2_4_BITS_102_TO_101_5_EQ_0_6_ETC___d85 :2'd0; 
  assign  RTL__IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137 =( RTL__stage2_rg_stage2 [100:96]==5'd0) ? 2'd0:(( RTL__near_mem$dmem_valid &&! RTL__near_mem$dmem_exc ) ? 2'd2:2'd1); 
  assign  RTL__IF_stage2_rg_stage2_4_BITS_102_TO_101_5_EQ_0_6_ETC___d85 =( RTL__stage2_rg_stage2 [102:101]==2'd0) ? 2'd2:( RTL__near_mem$dmem_valid  ? ( RTL__near_mem$dmem_exc  ? 2'd3:2'd2):2'd1); 
  assign  RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 = RTL__cur_verbosity__h1827 >4'd1; 
  assign  RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d730 = RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 &&( RTL__stage2_rg_stage2 [102:101]==2'd0|| RTL__near_mem$dmem_valid &&! RTL__near_mem$dmem_exc ); 
  assign  RTL__NOT_IF_stage2_rg_full_3_THEN_IF_stage2_rg_stag_ETC___d109 = RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3&&( RTL__stage2_rg_stage2 [102:101]==2'd0|| RTL__near_mem$dmem_valid &&! RTL__near_mem$dmem_exc ); 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 =! RTL__csr_regfile$interrupt_pending [4]&&! RTL__csr_regfile$nmi_pending ||(! RTL__stage1_rg_full || RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 )&&(! RTL__stage1_rg_full || RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 ); 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 =! RTL__csr_regfile$interrupt_pending [4]&&! RTL__csr_regfile$nmi_pending || RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 = RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 &&( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)&& RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ; 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 = RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 &&( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)&& RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ||! RTL__stage1_rg_full ; 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d769 =(! RTL__csr_regfile$interrupt_pending [4]&&! RTL__csr_regfile$nmi_pending || RTL___0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 )&& RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ; 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 =(! RTL__csr_regfile$interrupt_pending [4]&&! RTL__csr_regfile$nmi_pending || RTL___0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 )&&( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0); 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d776 = RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 &&( RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ||! RTL__stage1_rg_full ); 
  assign  RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d790 =! RTL__csr_regfile$interrupt_pending [4]&&! RTL__csr_regfile$nmi_pending ||! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ); 
  assign  RTL__NOT_near_mem_imem_exc__78_13_AND_IF_near_mem_i_ETC___d481 =! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd0&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd1&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd2&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd3&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd4&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd5&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd6&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd7&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd8&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd9&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd10; 
  assign  RTL__NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252 =( RTL__near_mem$imem_instr [14:12]!=3'b0|| RTL__near_mem$imem_instr [6:0]==7'b0110011&& RTL__near_mem$imem_instr [30])&&( RTL__near_mem$imem_instr [14:12]!=3'b0|| RTL__near_mem$imem_instr [6:0]!=7'b0110011||! RTL__near_mem$imem_instr [30])&& RTL__near_mem$imem_instr [14:12]!=3'b010&& RTL__near_mem$imem_instr [14:12]!=3'b011&& RTL__near_mem$imem_instr [14:12]!=3'b100&& RTL__near_mem$imem_instr [14:12]!=3'b110&& RTL__near_mem$imem_instr [14:12]!=3'b111; 
  assign  RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 =! RTL__near_mem$imem_valid || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd1&&( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 || RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 ); 
  assign  RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 = RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 ||! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ); 
  assign  RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 = RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 || RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL__SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 ={{20{ RTL__near_memimem_instr_BITS_31_TO_20__q7 [11]}}, RTL__near_memimem_instr_BITS_31_TO_20__q7 }; 
  assign  RTL___0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 = RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL___theResult_____1_fst__h6562 =( RTL__near_mem$imem_instr [14:12]==3'b0&& RTL__near_mem$imem_instr [6:0]==7'b0110011&& RTL__near_mem$imem_instr [30]) ?  RTL__rd_val___1__h6558 : RTL___theResult_____1_fst__h6569 ; 
  assign  RTL___theResult_____1_fst__h6597 = RTL__rs1_val_bypassed__h3337 & RTL___theResult___snd__h7382 ; 
  assign  RTL___theResult____h10743 =( RTL__delta_CPI_instrs__h10742 ==64'd0) ?  RTL__delta_CPI_instrs___1__h10778 : RTL__delta_CPI_instrs__h10742 ; 
  assign  RTL___theResult___snd__h7382 =( RTL__near_mem$imem_instr [6:0]==7'b0010011) ?  RTL__SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 : RTL__rs2_val__h5339 ; 
  assign  RTL__alu_outputs___1_addr__h5365 = RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  ?  RTL__alu_outputs___1_val2__h5367 : RTL__alu_outputs___1_val1__h5386 ; 
  assign  RTL__alu_outputs___1_addr__h5385 = RTL__near_mem$imem_pc +{{11{ RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 [20]}}, RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 }; 
  assign  RTL__alu_outputs___1_addr__h5410 ={ RTL__eaddr__h5553 [31:1],1'd0}; 
  assign  RTL__alu_outputs___1_addr__h5583 = RTL__rs1_val_bypassed__h3337 +{{20{ RTL__near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 [11]}}, RTL__near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 }; 
  assign  RTL__alu_outputs___1_exc_code__h5362 = RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616  ? 4'd0:4'd2; 
  assign  RTL__alu_outputs___1_exc_code__h5843 =( RTL__near_mem$imem_instr [14:12]==3'b0) ? (( RTL__near_mem$imem_instr [11:7]==5'd0&& RTL__near_mem$imem_instr [19:15]==5'd0) ?  RTL__CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4 :4'd2):4'd2; 
  assign  RTL__alu_outputs___1_val1__h5386 = RTL__near_mem$imem_pc +32'd4; 
  assign  RTL__alu_outputs___1_val1__h5480 =( RTL__near_mem$imem_instr [14:12]==3'b001) ?  RTL__rd_val__h7278 :( RTL__near_mem$imem_instr [30] ?  RTL__rd_val__h7352 : RTL__rd_val__h7330 ); 
  assign  RTL__alu_outputs___1_val1__h5516 =( RTL__near_mem$imem_instr [14:12]==3'b0&&( RTL__near_mem$imem_instr [6:0]!=7'b0110011||! RTL__near_mem$imem_instr [30])) ?  RTL__rd_val___1__h6550 : RTL___theResult_____1_fst__h6562 ; 
  assign  RTL__alu_outputs___1_val1__h5847 = RTL__near_mem$imem_instr [14] ? {27'd0, RTL__near_mem$imem_instr [19:15]}: RTL__rs1_val_bypassed__h3337 ; 
  assign  RTL__alu_outputs___1_val2__h5367 = RTL__near_mem$imem_pc +{{19{ RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 [12]}}, RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 }; 
  assign  RTL__cpi__h10745 = RTL__x__h10744 /64'd10; 
  assign  RTL__cpifrac__h10746 = RTL__x__h10744 %64'd10; 
  assign  RTL__csr_regfile_interrupt_pending_rg_cur_priv_9_07_ETC___d779 =( RTL__csr_regfile$interrupt_pending [4]|| RTL__csr_regfile$nmi_pending )&&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )|| RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd2&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0; 
  assign  RTL__csr_regfile_read_csr_mcycle__8_MINUS_rg_start__ETC___d818 = RTL__delta_CPI_cycles__h10741 *64'd10; 
  assign  RTL__cur_verbosity__h1827 =( RTL__csr_regfile$read_csr_minstret < RTL__cfg_logdelay ) ? 4'd0: RTL__cfg_verbosity ; 
  assign  RTL__data_to_stage2_addr__h5215 = RTL__x_out_data_to_stage2_addr__h5223 ; 
  assign  RTL__delta_CPI_cycles__h10741 = RTL__csr_regfile$read_csr_mcycle - RTL__rg_start_CPI_cycles ; 
  assign  RTL__delta_CPI_instrs___1__h10778 = RTL__delta_CPI_instrs__h10742 +64'd1; 
  assign  RTL__delta_CPI_instrs__h10742 = RTL__csr_regfile$read_csr_minstret - RTL__rg_start_CPI_instrs ; 
  assign  RTL__eaddr__h5553 = RTL__rs1_val_bypassed__h3337 + RTL__SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 ; 
  assign  RTL__fall_through_pc__h5175 = RTL__near_mem$imem_pc +( RTL__near_mem$imem_is_i32_not_i16  ? 32'd4:32'd2); 
  assign  RTL__gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 = RTL__gpr_regfile$RDY_server_reset_request_put && RTL__near_mem$RDY_server_reset_request_put && RTL__csr_regfile$RDY_server_reset_request_put && RTL__f_reset_reqs$EMPTY_N && RTL__stage1_f_reset_reqs$FULL_N && RTL__stage2_f_reset_reqs$FULL_N && RTL__stage3_f_reset_reqs$FULL_N ; 
  assign  RTL__gpr_regfile_RDY_server_reset_response_get__76__ETC___d688 = RTL__gpr_regfile$RDY_server_reset_response_get && RTL__near_mem$RDY_server_reset_response_get && RTL__csr_regfile$RDY_server_reset_response_get && RTL__stage1_f_reset_rsps$EMPTY_N && RTL__stage2_f_reset_rsps$EMPTY_N && RTL__stage3_f_reset_rsps$EMPTY_N && RTL__f_reset_rsps$FULL_N ; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d578 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd0; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d581 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd1; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d584 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd2; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d587 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd3; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d590 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd4; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d593 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd5; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d596 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd6; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d599 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd7; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d602 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd8; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d605 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd9; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d608 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd10; 
  assign  RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d611 =( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd0&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd1&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd2&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd3&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd4&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd5&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd6&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd7&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd8&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd9&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd10; 
  assign  RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328 = RTL__near_mem$imem_instr [14:12]==3'b0&&( RTL__near_mem$imem_instr [6:0]!=7'b0110011||! RTL__near_mem$imem_instr [30])|| RTL__near_mem$imem_instr [14:12]==3'b0&& RTL__near_mem$imem_instr [6:0]==7'b0110011&& RTL__near_mem$imem_instr [30]|| RTL__near_mem$imem_instr [14:12]==3'b010|| RTL__near_mem$imem_instr [14:12]==3'b011|| RTL__near_mem$imem_instr [14:12]==3'b100|| RTL__near_mem$imem_instr [14:12]==3'b110|| RTL__near_mem$imem_instr [14:12]==3'b111; 
  assign  RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616 =( RTL__near_mem$imem_instr [14:12]==3'b0|| RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b100|| RTL__near_mem$imem_instr [14:12]==3'b101|| RTL__near_mem$imem_instr [14:12]==3'b110|| RTL__near_mem$imem_instr [14:12]==3'b111)&& RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 && RTL__alu_outputs___1_val2__h5367 [1]; 
  assign  RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 = RTL__near_mem$imem_valid &&( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd1||! RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 &&! RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 ); 
  assign  RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 = RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&( RTL__near_mem$imem_exc || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ); 
  assign  RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 = RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ); 
  assign  RTL__near_memimem_instr_BITS_31_TO_20__q7 = RTL__near_mem$imem_instr [31:20]; 
  assign  RTL__near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 ={ RTL__near_mem$imem_instr [31:25], RTL__near_mem$imem_instr [11:7]}; 
  assign  RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 ={ RTL__near_mem$imem_instr [31], RTL__near_mem$imem_instr [7], RTL__near_mem$imem_instr [30:25], RTL__near_mem$imem_instr [11:8],1'b0}; 
  assign  RTL__near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 ={ RTL__near_mem$imem_instr [31], RTL__near_mem$imem_instr [19:12], RTL__near_mem$imem_instr [20], RTL__near_mem$imem_instr [30:21],1'b0}; 
  assign  RTL__output_stage2___1_bypass_rd_val__h4960 =(! RTL__near_mem$dmem_valid ||! RTL__near_mem$dmem_exc ) ? (( RTL__stage2_rg_stage2 [100:96]==5'd0) ?  RTL__stage2_rg_stage2 [63:32]: RTL__near_mem$dmem_word64 [31:0]): RTL__stage2_rg_stage2 [63:32]; 
  assign  RTL__rd_val___1__h6550 = RTL__rs1_val_bypassed__h3337 + RTL___theResult___snd__h7382 ; 
  assign  RTL__rd_val___1__h6558 = RTL__rs1_val_bypassed__h3337 - RTL___theResult___snd__h7382 ; 
  assign  RTL__rd_val___1__h6565 =(( RTL__rs1_val_bypassed__h3337 ^32'h80000000)<( RTL___theResult___snd__h7382 ^32'h80000000)) ? 32'd1:32'd0; 
  assign  RTL__rd_val___1__h6572 =( RTL__rs1_val_bypassed__h3337 < RTL___theResult___snd__h7382 ) ? 32'd1:32'd0; 
  assign  RTL__rd_val___1__h6579 = RTL__rs1_val_bypassed__h3337 ^ RTL___theResult___snd__h7382 ; 
  assign  RTL__rd_val___1__h6586 = RTL__rs1_val_bypassed__h3337 | RTL___theResult___snd__h7382 ; 
  assign  RTL__rd_val__h5072 =( RTL__stage3_rg_full && RTL__stage3_rg_stage3 [37]&& RTL__stage3_rg_stage3 [36:32]== RTL__near_mem$imem_instr [19:15]) ?  RTL__stage3_rg_stage3 [31:0]: RTL__gpr_regfile$read_rs1 ; 
  assign  RTL__rd_val__h5132 =( RTL__stage3_rg_full && RTL__stage3_rg_stage3 [37]&& RTL__stage3_rg_stage3 [36:32]== RTL__near_mem$imem_instr [24:20]) ?  RTL__stage3_rg_stage3 [31:0]: RTL__gpr_regfile$read_rs2 ; 
  assign  RTL__rd_val__h5523 ={ RTL__near_mem$imem_instr [31:12],12'h0}; 
  assign  RTL__rd_val__h5537 = RTL__near_mem$imem_pc + RTL__rd_val__h5523 ; 
  assign  RTL__rd_val__h7278 = RTL__rs1_val_bypassed__h3337 << RTL__shamt__h5467 ; 
  assign  RTL__rd_val__h7330 = RTL__rs1_val_bypassed__h3337 >> RTL__shamt__h5467 ; 
  assign  RTL__rd_val__h7352 = RTL__rs1_val_bypassed__h3337 >> RTL__shamt__h5467 |~(32'hFFFFFFFF>> RTL__shamt__h5467 )&{32{ RTL__rs1_val_bypassed__h3337 [31]}}; 
  assign  RTL__rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_EQ_0_ETC___d392 =( RTL__rg_cur_priv ==2'b11|| RTL__rg_cur_priv ==2'b01&&! RTL__csr_regfile$read_mstatus [21]|| RTL__rg_cur_priv ==2'b0&& RTL__csr_regfile$read_misa [13])&& RTL__near_mem$imem_instr [31:20]==12'b000100000101; 
  assign  RTL__rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 = RTL__rg_state ==4'd3&& RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d790 &&! RTL__stage3_rg_full && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0; 
  assign  RTL__rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 = RTL__rg_trap_info [67:36]== RTL__csr_regfile$csr_trap_actions [97:66]; 
  assign  RTL__rs1_val__h11213 =( RTL__rg_trap_instr [14:12]==3'b001) ?  RTL__rg_csr_val1 :{27'd0, RTL__rg_trap_instr [19:15]}; 
  assign  RTL__rs1_val_bypassed__h3337 =( RTL__near_mem$imem_instr [19:15]==5'd0) ? 32'd0: RTL__val__h5074 ; 
  assign  RTL__rs2_val__h5339 =( RTL__near_mem$imem_instr [24:20]==5'd0) ? 32'd0: RTL__val__h5134 ; 
  assign  RTL__shamt__h5467 =( RTL__near_mem$imem_instr [6:0]==7'b0010011) ?  RTL__near_mem$imem_instr [24:20]: RTL__rs2_val__h5339 [4:0]; 
  assign  RTL__trap_info_tval__h6925 = RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d649  ?  RTL__near_mem$imem_instr : RTL__IF_IF_near_mem_imem_instr__59_BITS_6_TO_0_79_E_ETC___d655 ; 
  assign  RTL__val__h5074 =( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd2&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 ) ?  RTL__x_out_bypass_rd_val__h4969 : RTL__rd_val__h5072 ; 
  assign  RTL__val__h5134 =( RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd2&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 ) ?  RTL__x_out_bypass_rd_val__h4969 : RTL__rd_val__h5132 ; 
  assign  RTL__value__h6967 = RTL__near_mem$imem_exc  ?  RTL__near_mem$imem_tval : RTL__trap_info_tval__h6925 ; 
  assign  RTL__x__h10744 = RTL__csr_regfile_read_csr_mcycle__8_MINUS_rg_start__ETC___d818 [63:0]/ RTL___theResult____h10743 ; 
  assign  RTL__x_exc_code__h15410 =( RTL__csr_regfile$interrupt_pending [4]&&! RTL__csr_regfile$nmi_pending ) ?  RTL__csr_regfile$interrupt_pending [3:0]:4'd0; 
  assign  RTL__x_out_bypass_rd_val__h4969 =( RTL__stage2_rg_stage2 [102:101]==2'd0) ?  RTL__stage2_rg_stage2 [63:32]: RTL__output_stage2___1_bypass_rd_val__h4960 ; 
  assign  RTL__x_out_data_to_stage2_rd__h5222 =( RTL__near_mem$imem_instr [6:0]==7'b1100011) ? 5'd0: RTL__near_mem$imem_instr [11:7]; 
  assign  RTL__x_out_data_to_stage2_val2__h5225 =( RTL__near_mem$imem_instr [6:0]==7'b1100011) ?  RTL__alu_outputs___1_val2__h5367 : RTL__rs2_val__h5339 ; 
  assign  RTL__x_out_next_pc__h5189 = RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  ?  RTL__data_to_stage2_addr__h5215 : RTL__fall_through_pc__h5175 ; 
  assign  RTL__x_out_trap_info_exc_code__h6928 = RTL__near_mem$imem_exc  ?  RTL__near_mem$imem_exc_code : RTL__alu_outputs_exc_code__h5862 ; 
  assign  RTL__y__h12191 =~ RTL__rs1_val__h11920 ; 
  always @(  RTL__stage2_rg_stage2  )
         begin 
             case ( RTL__stage2_rg_stage2 [102:101])
              2 'd0,2'd1: 
                  RTL__x_out_data_to_stage3_rd__h4667  = RTL__stage2_rg_stage2 [100:96];
              default : 
                  RTL__x_out_data_to_stage3_rd__h4667  =5'd0;endcase
         end
  always @(   RTL__stage2_rg_stage2            or   RTL__near_mem$dmem_word64  )
         begin 
             case ( RTL__stage2_rg_stage2 [102:101])
              2 'd0: 
                  RTL__x_out_data_to_stage3_rd_val__h4668  = RTL__stage2_rg_stage2 [63:32];
              2 'd1: 
                  RTL__x_out_data_to_stage3_rd_val__h4668  = RTL__near_mem$dmem_word64 [31:0];
              default : 
                  RTL__x_out_data_to_stage3_rd_val__h4668  = RTL__stage2_rg_stage2 [63:32];endcase
         end
  always @(   RTL__rg_trap_instr            or   RTL__rg_csr_val1  )
         begin 
             case ( RTL__rg_trap_instr [14:12])
              3 'b010,3'b011: 
                  RTL__rs1_val__h11920  = RTL__rg_csr_val1 ;
              default : 
                  RTL__rs1_val__h11920  ={27'd0, RTL__rg_trap_instr [19:15]};endcase
         end
  always @(  RTL__rg_cur_priv  )
         begin 
             case ( RTL__rg_cur_priv )
              2 'b0: 
                  RTL__CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  =4'd8;
              2 'b01: 
                  RTL__CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  =4'd9;
              default : 
                  RTL__CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  =4'd11;endcase
         end
  always @(   RTL__near_mem$imem_instr            or   RTL__CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  )
         begin 
             case ( RTL__near_mem$imem_instr [31:20])
              12 'b0: 
                  RTL__CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4  = RTL__CASE_rg_cur_priv_0b0_8_0b1_9_11__q3 ;
              12 'b000000000001: 
                  RTL__CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4  =4'd3;
              default : 
                  RTL__CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4  =4'd2;endcase
         end
  always @(     RTL__stage2_rg_stage2                or   RTL__near_mem$dmem_valid            or   RTL__near_mem$dmem_exc           or   RTL__IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137  )
         begin 
             case ( RTL__stage2_rg_stage2 [102:101])
              2 'd0: 
                  RTL__CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5  =2'd2;
              2 'd1: 
                  RTL__CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5  =(! RTL__near_mem$dmem_valid ||! RTL__near_mem$dmem_exc ) ?  RTL__IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137 :2'd0;
              default : 
                  RTL__CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5  =2'd0;endcase
         end
  always @(     RTL__near_mem$imem_instr                or   RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220            or   RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216           or   RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b001: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  =! RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b100: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b101: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  =! RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b110: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL__near_mem$imem_instr [14:12]==3'b111&&! RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;endcase
         end
  always @(       RTL__near_mem$imem_instr                    or   RTL__alu_outputs___1_addr__h5583              or   RTL__eaddr__h5553             or   RTL__alu_outputs___1_addr__h5365            or   RTL__alu_outputs___1_addr__h5410           or   RTL__alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0000011: 
                  RTL__x_out_data_to_stage2_addr__h5223  = RTL__eaddr__h5553 ;
              7 'b1100011: 
                  RTL__x_out_data_to_stage2_addr__h5223  = RTL__alu_outputs___1_addr__h5365 ;
              7 'b1100111: 
                  RTL__x_out_data_to_stage2_addr__h5223  = RTL__alu_outputs___1_addr__h5410 ;
              7 'b1101111: 
                  RTL__x_out_data_to_stage2_addr__h5223  = RTL__alu_outputs___1_addr__h5385 ;
              default : 
                  RTL__x_out_data_to_stage2_addr__h5223  = RTL__alu_outputs___1_addr__h5583 ;endcase
         end
  always @(       RTL__near_mem$imem_instr                    or   RTL___theResult_____1_fst__h6597              or   RTL__rd_val___1__h6565             or   RTL__rd_val___1__h6572            or   RTL__rd_val___1__h6579           or   RTL__rd_val___1__h6586  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b010: 
                  RTL___theResult_____1_fst__h6569  = RTL__rd_val___1__h6565 ;
              3 'b011: 
                  RTL___theResult_____1_fst__h6569  = RTL__rd_val___1__h6572 ;
              3 'b100: 
                  RTL___theResult_____1_fst__h6569  = RTL__rd_val___1__h6579 ;
              3 'b110: 
                  RTL___theResult_____1_fst__h6569  = RTL__rd_val___1__h6586 ;
              default : 
                  RTL___theResult_____1_fst__h6569  = RTL___theResult_____1_fst__h6597 ;endcase
         end
  always @(     RTL__near_mem$imem_instr                or   RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220            or   RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216           or   RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  =! RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b001: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  = RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b100: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  =! RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b101: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  = RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b110: 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  =! RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  = RTL__near_mem$imem_instr [14:12]!=3'b111|| RTL__IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;endcase
         end
  always @(   RTL__near_mem$imem_instr            or   RTL__NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0010011,7'b0110011: 
                  RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8  = RTL__NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252 ;
              default : 
                  RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8  = RTL__near_mem$imem_instr [6:0]!=7'b0110111&& RTL__near_mem$imem_instr [6:0]!=7'b0010111&&(( RTL__near_mem$imem_instr [6:0]==7'b0000011) ?  RTL__near_mem$imem_instr [14:12]!=3'b0&& RTL__near_mem$imem_instr [14:12]!=3'b100&& RTL__near_mem$imem_instr [14:12]!=3'b001&& RTL__near_mem$imem_instr [14:12]!=3'b101&& RTL__near_mem$imem_instr [14:12]!=3'b010: RTL__near_mem$imem_instr [6:0]!=7'b0100011|| RTL__near_mem$imem_instr [14:12]!=3'b0&& RTL__near_mem$imem_instr [14:12]!=3'b001&& RTL__near_mem$imem_instr [14:12]!=3'b010);endcase
         end
  always @(      RTL__near_mem$imem_instr                  or   RTL__eaddr__h5553             or   RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285            or   RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291           or   RTL__alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b1100011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308  = RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285 || RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 ;
              7 'b1101111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308  = RTL__alu_outputs___1_addr__h5385 [1];
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308  = RTL__near_mem$imem_instr [6:0]!=7'b1100111|| RTL__eaddr__h5553 [1];endcase
         end
  always @(   RTL__near_mem$imem_instr            or   RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0010011,7'b0110011: 
                  RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9  = RTL__near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328 ;
              default : 
                  RTL__CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9  = RTL__near_mem$imem_instr [6:0]==7'b0110111|| RTL__near_mem$imem_instr [6:0]==7'b0010111||(( RTL__near_mem$imem_instr [6:0]==7'b0000011) ?  RTL__near_mem$imem_instr [14:12]==3'b0|| RTL__near_mem$imem_instr [14:12]==3'b100|| RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b101|| RTL__near_mem$imem_instr [14:12]==3'b010: RTL__near_mem$imem_instr [6:0]==7'b0100011&&( RTL__near_mem$imem_instr [14:12]==3'b0|| RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b010));endcase
         end
  always @(       RTL__near_mem$imem_instr                    or   RTL__eaddr__h5553              or   RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291             or   RTL__alu_outputs___1_val2__h5367            or   RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227           or   RTL__alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b1100011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  =( RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 ||! RTL__alu_outputs___1_val2__h5367 [1])&&( RTL__near_mem$imem_instr [14:12]==3'b0|| RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b100|| RTL__near_mem$imem_instr [14:12]==3'b101|| RTL__near_mem$imem_instr [14:12]==3'b110|| RTL__near_mem$imem_instr [14:12]==3'b111)&& RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 ;
              7 'b1101111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  =! RTL__alu_outputs___1_addr__h5385 [1];
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  = RTL__near_mem$imem_instr [6:0]==7'b1100111&&! RTL__eaddr__h5553 [1];endcase
         end
  always @(    RTL__near_mem$imem_instr              or   RTL__rg_cur_priv           or   RTL__IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394  )
         begin 
             case ( RTL__near_mem$imem_instr [31:20])
              12 'b0,12'b000000000001: 
                  RTL__IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396  =4'd11;
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396  =( RTL__rg_cur_priv ==2'b11&& RTL__near_mem$imem_instr [31:20]==12'b001100000010) ? 4'd7: RTL__IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394 ;endcase
         end
  always @(  RTL__near_mem$imem_instr  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b0,3'b001,3'b010,3'b100,3'b101: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10  =4'd0;
              default : 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10  =4'd11;endcase
         end
  always @(  RTL__near_mem$imem_instr  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11  =4'd4;
              3 'b001: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11  =4'd5;
              default : 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11  =4'd11;endcase
         end
  always @(  RTL__near_mem$imem_instr  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b0,3'b001,3'b010: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12  =4'd0;
              default : 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12  =4'd11;endcase
         end
  always @(   RTL__near_mem$imem_instr            or   RTL__IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396  )
         begin 
             case ( RTL__near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =( RTL__near_mem$imem_instr [11:7]==5'd0&& RTL__near_mem$imem_instr [19:15]==5'd0) ?  RTL__IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396 :4'd11;
              3 'b001,3'b101: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =4'd2;
              3 'b010,3'b011,3'b110,3'b111: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =4'd3;
              3 'd4: 
                  RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =4'd11;endcase
         end
  always @(       RTL__near_mem$imem_instr                    or   RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10              or   RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11             or   RTL__IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362            or   RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12           or   RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0000011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10 ;
              7 'b0001111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11 ;
              7 'b0010011,7'b0110011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL__IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362 ;
              7 'b0010111,7'b0110111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  =4'd0;
              7 'b0100011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12 ;
              7 'b1110011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL__CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13 ;
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  =4'd11;endcase
         end
  always @(       RTL__near_mem$imem_instr                    or   RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409              or   RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285             or   RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227            or   RTL__eaddr__h5553           or   RTL__alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b1100011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  = RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285  ? 4'd11:( RTL__IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  ? 4'd1:4'd0);
              7 'b1100111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  = RTL__eaddr__h5553 [1] ? 4'd11:4'd1;
              7 'b1101111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  = RTL__alu_outputs___1_addr__h5385 [1] ? 4'd11:4'd1;
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  =(( RTL__near_mem$imem_instr [6:0]==7'b0010011|| RTL__near_mem$imem_instr [6:0]==7'b0110011)&&( RTL__near_mem$imem_instr [14:12]==3'b001|| RTL__near_mem$imem_instr [14:12]==3'b101)) ? ( RTL__near_mem$imem_instr [25] ? 4'd11:4'd0): RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409 ;endcase
         end
  always @(  RTL__near_mem$imem_instr  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0000011: 
                  RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491  =2'd1;
              7 'b0010011,7'b0010111,7'b0110011,7'b0110111,7'b1100011,7'b1100111,7'b1101111: 
                  RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491  =2'd0;
              default : 
                  RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491  =2'd2;endcase
         end
  always @(    RTL__near_mem$imem_instr              or   RTL__alu_outputs___1_exc_code__h5362           or   RTL__alu_outputs___1_exc_code__h5843  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0000011,7'b0001111,7'b0010011,7'b0010111,7'b0100011,7'b0110011,7'b0110111: 
                  RTL__alu_outputs_exc_code__h5862  =4'd2;
              7 'b1100011: 
                  RTL__alu_outputs_exc_code__h5862  = RTL__alu_outputs___1_exc_code__h5362 ;
              7 'b1100111,7'b1101111: 
                  RTL__alu_outputs_exc_code__h5862  =4'd0;
              7 'b1110011: 
                  RTL__alu_outputs_exc_code__h5862  = RTL__alu_outputs___1_exc_code__h5843 ;
              default : 
                  RTL__alu_outputs_exc_code__h5862  =4'd2;endcase
         end
  always @(      RTL__near_mem$imem_instr                  or   RTL__alu_outputs___1_val1__h5847             or   RTL__alu_outputs___1_val1__h5516            or   RTL__rd_val__h5537           or   RTL__rd_val__h5523  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b0010011,7'b0110011: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL__alu_outputs___1_val1__h5516 ;
              7 'b0010111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL__rd_val__h5537 ;
              7 'b0110111: 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL__rd_val__h5523 ;
              default : 
                  RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL__alu_outputs___1_val1__h5847 ;endcase
         end
  always @(    RTL__near_mem$imem_instr              or   RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571           or   RTL__alu_outputs___1_val1__h5386  )
         begin 
             case ( RTL__near_mem$imem_instr [6:0])
              7 'b1100111,7'b1101111: 
                  RTL__x_out_data_to_stage2_val1__h5224  = RTL__alu_outputs___1_val1__h5386 ;
              default : 
                  RTL__x_out_data_to_stage2_val1__h5224  = RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571 ;endcase
         end
  always @( posedge  RTL__CLK )
         begin 
             if ( RTL__RST_N ==1'b0)
                 begin  
                     RTL__cfg_logdelay  <=64'd0; 
                     RTL__cfg_verbosity  <=4'd0; 
                     RTL__rg_cur_priv  <=2'b11; 
                     RTL__rg_retiring  <=1'd0; 
                     RTL__rg_run_on_reset  <=1'd0; 
                     RTL__rg_state  <=4'd0; 
                     RTL__s1_to_s2  <=1'd0; 
                     RTL__s2_to_s3  <=1'd0; 
                     RTL__s3_deq  <=1'd0; 
                     RTL__stage1_rg_full  <=1'd0; 
                     RTL__stage2_rg_full  <=1'd0; 
                     RTL__stage2_rg_resetting  <=1'd0; 
                     RTL__stage3_rg_full  <=1'd0;
                 end 
              else 
                 begin 
                     if ( RTL__cfg_logdelay$EN ) 
                         RTL__cfg_logdelay  <= RTL__cfg_logdelay$D_IN ;
                     if ( RTL__cfg_verbosity$EN ) 
                         RTL__cfg_verbosity  <= RTL__cfg_verbosity$D_IN ;
                     if ( RTL__rg_cur_priv$EN ) 
                         RTL__rg_cur_priv  <= RTL__rg_cur_priv$D_IN ;
                     if ( RTL__rg_retiring$EN ) 
                         RTL__rg_retiring  <= RTL__rg_retiring$D_IN ;
                     if ( RTL__rg_run_on_reset$EN ) 
                         RTL__rg_run_on_reset  <= RTL__rg_run_on_reset$D_IN ;
                     if ( RTL__rg_state$EN ) 
                         RTL__rg_state  <= RTL__rg_state$D_IN ;
                     if ( RTL__s1_to_s2$EN ) 
                         RTL__s1_to_s2  <= RTL__s1_to_s2$D_IN ;
                     if ( RTL__s2_to_s3$EN ) 
                         RTL__s2_to_s3  <= RTL__s2_to_s3$D_IN ;
                     if ( RTL__s3_deq$EN ) 
                         RTL__s3_deq  <= RTL__s3_deq$D_IN ;
                     if ( RTL__stage1_rg_full$EN ) 
                         RTL__stage1_rg_full  <= RTL__stage1_rg_full$D_IN ;
                     if ( RTL__stage2_rg_full$EN ) 
                         RTL__stage2_rg_full  <= RTL__stage2_rg_full$D_IN ;
                     if ( RTL__stage2_rg_resetting$EN ) 
                         RTL__stage2_rg_resetting  <= RTL__stage2_rg_resetting$D_IN ;
                     if ( RTL__stage3_rg_full$EN ) 
                         RTL__stage3_rg_full  <= RTL__stage3_rg_full$D_IN ;
                 end 
             if ( RTL__rg_csr_pc$EN ) 
                 RTL__rg_csr_pc  <= RTL__rg_csr_pc$D_IN ;
             if ( RTL__rg_csr_val1$EN ) 
                 RTL__rg_csr_val1  <= RTL__rg_csr_val1$D_IN ;
             if ( RTL__rg_mstatus_MXR$EN ) 
                 RTL__rg_mstatus_MXR  <= RTL__rg_mstatus_MXR$D_IN ;
             if ( RTL__rg_next_pc$EN ) 
                 RTL__rg_next_pc  <= RTL__rg_next_pc$D_IN ;
             if ( RTL__rg_sstatus_SUM$EN ) 
                 RTL__rg_sstatus_SUM  <= RTL__rg_sstatus_SUM$D_IN ;
             if ( RTL__rg_start_CPI_cycles$EN ) 
                 RTL__rg_start_CPI_cycles  <= RTL__rg_start_CPI_cycles$D_IN ;
             if ( RTL__rg_start_CPI_instrs$EN ) 
                 RTL__rg_start_CPI_instrs  <= RTL__rg_start_CPI_instrs$D_IN ;
             if ( RTL__rg_trap_info$EN ) 
                 RTL__rg_trap_info  <= RTL__rg_trap_info$D_IN ;
             if ( RTL__rg_trap_instr$EN ) 
                 RTL__rg_trap_instr  <= RTL__rg_trap_instr$D_IN ;
             if ( RTL__rg_trap_interrupt$EN ) 
                 RTL__rg_trap_interrupt  <= RTL__rg_trap_interrupt$D_IN ;
             if ( RTL__stage2_rg_stage2$EN ) 
                 RTL__stage2_rg_stage2  <= RTL__stage2_rg_stage2$D_IN ;
             if ( RTL__stage3_rg_stage3$EN ) 
                 RTL__stage3_rg_stage3  <= RTL__stage3_rg_stage3$D_IN ;
         end
  always @( negedge  RTL__CLK )
         begin #0;
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$display("================================================================");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$display("%0d: Pipeline State:  minstret:%0d  cur_priv:%0d  mstatus:%0x", RTL__csr_regfile$read_csr_mcycle , RTL__csr_regfile$read_csr_minstret , RTL__rg_cur_priv , RTL__csr_regfile$read_mstatus );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("    ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("MStatus{","sd:%0d", RTL__csr_regfile$read_mstatus [14:13]==2'h3|| RTL__csr_regfile$read_mstatus [16:15]==2'h3);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__csr_regfile$read_misa [27:26]==2'd2)$write(" sxl:%0d uxl:%0d",2'd0,2'd0);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__csr_regfile$read_misa [27:26]!=2'd2)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" tsr:%0d", RTL__csr_regfile$read_mstatus [22]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" tw:%0d", RTL__csr_regfile$read_mstatus [21]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" tvm:%0d", RTL__csr_regfile$read_mstatus [20]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" mxr:%0d", RTL__csr_regfile$read_mstatus [19]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" sum:%0d", RTL__csr_regfile$read_mstatus [18]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" mprv:%0d", RTL__csr_regfile$read_mstatus [17]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" xs:%0d", RTL__csr_regfile$read_mstatus [16:15]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" fs:%0d", RTL__csr_regfile$read_mstatus [14:13]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" mpp:%0d", RTL__csr_regfile$read_mstatus [12:11]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" spp:%0d", RTL__csr_regfile$read_mstatus [8]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" pies:%0d_%0d%0d", RTL__csr_regfile$read_mstatus [7], RTL__csr_regfile$read_mstatus [5], RTL__csr_regfile$read_mstatus [4]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write(" ies:%0d_%0d%0d", RTL__csr_regfile$read_mstatus [3], RTL__csr_regfile$read_mstatus [1], RTL__csr_regfile$read_mstatus [0]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("}");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("    Stage3: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("Output_Stage3");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage3_rg_full )$write(" PIPE");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage3_rg_full )$write(" EMPTY");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("        Bypass  to Stage1: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("Bypass {");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&(! RTL__stage3_rg_full ||! RTL__stage3_rg_stage3 [37]))$write("Rd -");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage3_rg_full && RTL__stage3_rg_stage3 [37])$write("Rd %0d ", RTL__stage3_rg_stage3 [36:32],"rd_val:%h", RTL__stage3_rg_stage3 [31:0]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("}");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$display("    Stage2: pc 0x%08h instr 0x%08h priv %0d", RTL__stage2_rg_stage2 [166:135], RTL__stage2_rg_stage2 [134:103], RTL__stage2_rg_stage2 [168:167]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("        ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("Output_Stage2"," EMPTY");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("Output_Stage2"," BUSY: pc:%0h", RTL__stage2_rg_stage2 [166:135]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("Output_Stage2"," NONPIPE: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("Output_Stage2"," PIPE: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("data_to_Stage3 {pc:%h  instr:%h  priv:%0d\n", RTL__stage2_rg_stage2 [166:135], RTL__stage2_rg_stage2 [134:103], RTL__stage2_rg_stage2 [168:167]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("        rd_valid:");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3&& RTL__stage2_rg_stage2 [102:101]!=2'd0&&(! RTL__near_mem$dmem_valid || RTL__near_mem$dmem_exc ))$write("False");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__NOT_IF_stage2_rg_full_3_THEN_IF_stage2_rg_stag_ETC___d109 )$write("True");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("  grd:%0d  rd_val:%h\n", RTL__x_out_data_to_stage3_rd__h4667 , RTL__x_out_data_to_stage3_rd_val__h4668 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("Trap_Info { ","epc: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL__stage2_rg_stage2 [166:135]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","exc_code: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL__near_mem$dmem_exc_code );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","tval: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL__stage2_rg_stage2 [95:64]," }");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(" ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("Trap_Info { ","epc: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL__stage2_rg_stage2 [166:135]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","exc_code: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL__near_mem$dmem_exc_code );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","tval: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL__stage2_rg_stage2 [95:64]," }");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("        Bypass  to Stage1: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("Bypass {");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd0)$write("Rd -");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd0)$write("Rd %0d ", RTL__stage2_rg_stage2 [100:96]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd0)$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd1)$write("-");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd0&& RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd1)$write("rd_val:%h", RTL__x_out_bypass_rd_val__h4969 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("}");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$display("    Stage1: pc 0x%08h instr 0x%08h priv %0d", RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("        ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("Output_Stage1"," BUSY pc:%h", RTL__near_mem$imem_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("Output_Stage1"," NONPIPE: pc:%h", RTL__near_mem$imem_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("Output_Stage1");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("Output_Stage1"," EMPTY");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write(" PIPE: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd0)$write("CONTROL_STRAIGHT");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd1)$write("CONTROL_BRANCH");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd2)$write("CONTROL_CSRR_W");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd3)$write("CONTROL_CSRR_S_or_C");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd4)$write("CONTROL_FENCE");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd5)$write("CONTROL_FENCE_I");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd6)$write("CONTROL_SFENCE_VMA");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd7)$write("CONTROL_MRET");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd8)$write("CONTROL_SRET");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd9)$write("CONTROL_URET");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd10)$write("CONTROL_WFI");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__NOT_near_mem_imem_exc__78_13_AND_IF_near_mem_i_ETC___d481 )$write("CONTROL_TRAP");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write(" ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("}");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("data_to_Stage 2 {pc:%h  instr:%h  priv:%0d\n", RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("            op_stage2:");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd0)$write("OP_Stage2_ALU");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd1)$write("OP_Stage2_LD");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL__near_mem$imem_exc &&( RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL__IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd0&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd1)$write("OP_Stage2_ST");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("  rd:%0d\n", RTL__x_out_data_to_stage2_rd__h5222 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("            addr:%h  val1:%h  val2:%h}", RTL__x_out_data_to_stage2_addr__h5223 , RTL__x_out_data_to_stage2_val1__h5224 , RTL__x_out_data_to_stage2_val2__h5225 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(" ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d578 )$write("CONTROL_STRAIGHT");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d581 )$write("CONTROL_BRANCH");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d584 )$write("CONTROL_CSRR_W");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d587 )$write("CONTROL_CSRR_S_or_C");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d590 )$write("CONTROL_FENCE");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d593 )$write("CONTROL_FENCE_I");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d596 )$write("CONTROL_SFENCE_VMA");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d599 )$write("CONTROL_MRET");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d602 )$write("CONTROL_SRET");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d605 )$write("CONTROL_URET");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d608 )$write("CONTROL_WFI");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL__near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d611 )$write("CONTROL_TRAP");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(" ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("Trap_Info { ","epc: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("'h%h", RTL__near_mem$imem_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(", ","exc_code: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("'h%h", RTL__x_out_trap_info_exc_code__h6928 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(", ","tval: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("'h%h", RTL__value__h6967 ," }");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe && RTL__stage1_rg_full && RTL__NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe &&! RTL__stage1_rg_full )$write("");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_show_pipe )$display("----------------");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__soc_map$m_pc_reset_value [31:0]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_complete && RTL__rg_run_on_reset )$display("%0d: %m.rl_reset_complete: restart at PC = 0x%0h", RTL__csr_regfile$read_csr_mcycle , RTL__soc_map$m_pc_reset_value [31:0]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_complete &&! RTL__rg_run_on_reset )$display("%0d: %m.rl_reset_complete: entering DEBUG_MODE", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_pipe", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__stage3_rg_full && RTL__stage3_rg_stage3 [37]&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    S3.fa_deq: write GRd 0x%0h, rd_val 0x%0h", RTL__stage3_rg_stage3 [36:32], RTL__stage3_rg_stage3 [31:0]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("    S3.enq: ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("data_to_Stage3 {pc:%h  instr:%h  priv:%0d\n", RTL__stage2_rg_stage2 [166:135], RTL__stage2_rg_stage2 [134:103], RTL__stage2_rg_stage2 [168:167]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("        rd_valid:");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL__stage2_rg_stage2 [102:101]!=2'd0&&(! RTL__near_mem$dmem_valid || RTL__near_mem$dmem_exc ))$write("False");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d730 )$write("True");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("  grd:%0d  rd_val:%h\n", RTL__x_out_data_to_stage3_rd__h4667 , RTL__x_out_data_to_stage3_rd_val__h4668 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__stage2_rg_stage2 [166:135], RTL__stage2_rg_stage2 [134:103], RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("    CPU_Stage2.enq (Data_Stage1_to_Stage2) ");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("data_to_Stage 2 {pc:%h  instr:%h  priv:%0d\n", RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("            op_stage2:");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd0)$write("OP_Stage2_ALU");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd1)$write("OP_Stage2_LD");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd0&& RTL__IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd1)$write("OP_Stage2_ST");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("  rd:%0d\n", RTL__x_out_data_to_stage2_rd__h5222 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("            addr:%h  val1:%h  val2:%h}", RTL__x_out_data_to_stage2_addr__h5223 , RTL__x_out_data_to_stage2_val1__h5224 , RTL__x_out_data_to_stage2_val2__h5225 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("\n");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_pipe && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 && RTL__NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__x_out_next_pc__h5189 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage2_nonpipe && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage2_nonpipe", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_trap && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_trap", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_trap && RTL__rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 )$display("%0d: %m.rl_stage1_trap: Tight infinite trap loop: pc 0x%0x instr 0x%08x", RTL__csr_regfile$read_csr_mcycle , RTL__csr_regfile$csr_trap_actions [97:66], RTL__rg_trap_instr );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_trap && RTL__rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 )$display("CPI: %0d.%0d = (%0d/%0d) since last 'continue'", RTL__cpi__h10745 , RTL__cpifrac__h10746 , RTL__delta_CPI_cycles__h10741 , RTL___theResult____h10743 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_trap && RTL__rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 )$finish(32'd0);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_trap && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__rg_trap_info [67:36], RTL__rg_trap_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_trap && RTL__cur_verbosity__h1827 !=4'd0)$display("    mcause:0x%0h  epc 0x%0h  tval:0x%0h  next_pc 0x%0h, new_priv %0d new_mstatus 0x%0h", RTL__csr_regfile$csr_trap_actions [33:2], RTL__rg_trap_info [67:36], RTL__rg_trap_info [31:0], RTL__csr_regfile$csr_trap_actions [97:66], RTL__csr_regfile$csr_trap_actions [1:0], RTL__csr_regfile$csr_trap_actions [65:34]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_W && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_W", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_W_2", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__rg_csr_pc , RTL__rg_trap_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL__csr_regfile$access_permitted_1 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    S1: write CSRRW/CSRRWI Rs1 %0d Rs1_val 0x%0h csr 0x%0h csr_val 0x%0h Rd %0d", RTL__rg_trap_instr [19:15], RTL__rs1_val__h11213 , RTL__rg_trap_instr [31:20], RTL__csr_regfile$read_csr [31:0], RTL__rg_trap_instr [11:7]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_W_2 &&! RTL__csr_regfile$access_permitted_1 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    rl_stage1_CSRR_W: Trap on CSR permissions: Rs1 %0d Rs1_val 0x%0h csr 0x%0h Rd %0d", RTL__rg_trap_instr [19:15], RTL__rs1_val__h11213 , RTL__rg_trap_instr [31:20], RTL__rg_trap_instr [11:7]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_S_or_C", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_S_or_C_2", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__rg_csr_pc , RTL__rg_trap_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL__csr_regfile$access_permitted_2 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    S1: write CSRR_S_or_C: Rs1 %0d Rs1_val 0x%0h csr 0x%0h csr_val 0x%0h Rd %0d", RTL__rg_trap_instr [19:15], RTL__rs1_val__h11920 , RTL__rg_trap_instr [31:20], RTL__csr_regfile$read_csr [31:0], RTL__rg_trap_instr [11:7]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 &&! RTL__csr_regfile$access_permitted_2 && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    rl_stage1_CSRR_S_or_C: Trap on CSR permissions: Rs1 %0d Rs1_val 0x%0h csr 0x%0h Rd %0d", RTL__rg_trap_instr [19:15], RTL__rs1_val__h11920 , RTL__rg_trap_instr [31:20], RTL__rg_trap_instr [11:7]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__x_out_next_pc__h5189 );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_restart_after_csrrx && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: rl_stage1_restart_after_csrrx: minstret:%0d  pc:%0x  cur_priv:%0d", RTL__csr_regfile$read_csr_mcycle , RTL__csr_regfile$read_csr_minstret , RTL__x_out_next_pc__h5189 , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_xRET && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_xRET", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_xRET && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_xRET && RTL__cur_verbosity__h1827 !=4'd0)$display("    xRET: next_pc:0x%0h  new mstatus:0x%0h  new priv:%0d", RTL__csr_regfile$csr_ret_actions [65:34], RTL__csr_regfile$csr_ret_actions [31:0], RTL__csr_regfile$csr_ret_actions [33:32]);
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_FENCE_I && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE_I", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_FENCE_I && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_FENCE_I && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE_I", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_FENCE_I && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_finish_FENCE_I", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_FENCE_I && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__rg_next_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_FENCE_I && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_finish_FENCE_I");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_FENCE && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_FENCE && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_FENCE && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_FENCE && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_finish_FENCE", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_FENCE && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__rg_next_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_FENCE && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_finish_FENCE");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_SFENCE_VMA", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_SFENCE_VMA && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_SFENCE_VMA", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_finish_SFENCE_VMA", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__rg_next_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_finish_SFENCE_VMA && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_finish_SFENCE_VMA");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_WFI && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_WFI", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_WFI && RTL__cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL__csr_regfile$read_csr_minstret , RTL__near_mem$imem_pc , RTL__near_mem$imem_instr , RTL__rg_cur_priv );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_WFI && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_stage1_WFI");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_WFI_resume && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_WFI_resume", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_WFI_resume && RTL__cur_verbosity__h1827 !=4'd0)$display("    WFI resume");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_WFI_resume && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__rg_next_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_from_WFI && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_reset_from_WFI", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_trap_fetch && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL__rg_next_pc );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_stage1_interrupt && RTL__NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_interrupt", RTL__csr_regfile$read_csr_mcycle );
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_start )$display("================================================================");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_start )$write("CPU: Bluespec  RISC-V  Piccolo  v3.0");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_start )$display(" (RV32)");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_start )$display("Copyright (c) 2016-2019 Bluespec, Inc. All Rights Reserved.");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_start )$display("================================================================");
             if ( RTL__RST_N !=1'b0)
                 if ( RTL__WILL_FIRE_RL_rl_reset_start && RTL__cur_verbosity__h1827 !=4'd0)$display("%0d: %m.rl_reset_start", RTL__csr_regfile$read_csr_mcycle );
         end
  assign  RTL__RTL__DOT__s3_deq$D_IN = RTL__s3_deq$D_IN ; 
  assign  RTL__RTL__DOT__near_mem$dmem_exc = RTL__near_mem$dmem_exc ; 
  assign  RTL__RTL__DOT__near_mem$imem_pc = RTL__near_mem$imem_pc ; 
  assign  RTL__RTL__DOT__near_mem$imem_instr = RTL__near_mem$imem_instr ; 
  assign  RTL__RTL__DOT__near_mem$dmem_req_addr = RTL__near_mem$dmem_req_addr ; 
  assign  RTL__RTL__DOT__stage2_rg_stage2 = RTL__stage2_rg_stage2 ; 
  assign  RTL__RTL__DOT__rg_cur_priv = RTL__rg_cur_priv ; 
  assign  RTL__RTL__DOT__near_mem$EN_dmem_req = RTL__near_mem$EN_dmem_req ; 
  assign  RTL__RTL__DOT__near_mem$dmem_req_f3 = RTL__near_mem$dmem_req_f3 ; 
  assign  RTL__RTL__DOT__s1_to_s2$D_IN = RTL__s1_to_s2$D_IN ; 
  assign  RTL__RTL__DOT__near_mem$dmem_word64 = RTL__near_mem$dmem_word64 ; 
  assign  RTL__RTL__DOT__stage3_rg_full = RTL__stage3_rg_full ; 
  assign  RTL__RTL__DOT__rg_trap_instr = RTL__rg_trap_instr ; 
  assign  RTL__RTL__DOT__near_mem$dmem_req_op = RTL__near_mem$dmem_req_op ; 
  assign  RTL__RTL__DOT__s2_to_s3$D_IN = RTL__s2_to_s3$D_IN ; 
  assign  RTL__RTL__DOT__rg_retiring$EN = RTL__rg_retiring$EN ; 
  assign  RTL__RTL__DOT__rg_state = RTL__rg_state ; 
  assign  RTL__RTL__DOT__s3_deq$EN = RTL__s3_deq$EN ; 
  assign  RTL__RTL__DOT__s1_to_s2$EN = RTL__s1_to_s2$EN ; 
  assign  RTL__RTL__DOT__s2_to_s3$EN = RTL__s2_to_s3$EN ; 
  assign  RTL__RTL__DOT__rg_run_on_reset = RTL__rg_run_on_reset ; 
  assign  RTL__RTL__DOT__stage1_rg_full = RTL__stage1_rg_full ; 
  assign  RTL__RTL__DOT__stage2_rg_full = RTL__stage2_rg_full ; 
  assign  RTL__RTL__DOT__near_mem$dmem_req_store_value = RTL__near_mem$dmem_req_store_value ;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__DOT__near_mem$dmem_req_op = RTL__RTL__DOT__near_mem$dmem_req_op;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__rg_trap_instr = RTL__RTL__DOT__rg_trap_instr;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL__RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__near_mem$dmem_req_store_value = RTL__RTL__DOT__near_mem$dmem_req_store_value;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__DOT__near_mem$dmem_word64 = RTL__RTL__DOT__near_mem$dmem_word64;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL__RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__s1_to_s2$D_IN = RTL__RTL__DOT__s1_to_s2$D_IN;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    assign RTL__DOT__stage2_rg_full = RTL__RTL__DOT__stage2_rg_full;
    assign RTL__DOT__csr_regfile__DOT__rg_state = RTL__RTL__DOT__csr_regfile__DOT__rg_state;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__DOT__stage1_rg_full = RTL__RTL__DOT__stage1_rg_full;
    assign RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    assign RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL__RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__rg_run_on_reset = RTL__RTL__DOT__rg_run_on_reset;
    assign RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL__RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL__RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__s2_to_s3$EN = RTL__RTL__DOT__s2_to_s3$EN;
    assign RTL__DOT__near_mem$dmem_req_f3 = RTL__RTL__DOT__near_mem$dmem_req_f3;
    assign RTL__DOT__s1_to_s2$EN = RTL__RTL__DOT__s1_to_s2$EN;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    assign RTL__DOT__s3_deq$EN = RTL__RTL__DOT__s3_deq$EN;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__rg_state = RTL__RTL__DOT__rg_state;
    assign RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__rg_retiring$EN = RTL__RTL__DOT__rg_retiring$EN;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__DOT__s2_to_s3$D_IN = RTL__RTL__DOT__s2_to_s3$D_IN;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    assign RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__stage3_rg_full = RTL__RTL__DOT__stage3_rg_full;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    assign RTL__DOT__stage2_rg_stage2 = RTL__RTL__DOT__stage2_rg_stage2;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    assign RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__csr_regfile__DOT__rg_nmi = RTL__RTL__DOT__csr_regfile__DOT__rg_nmi;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL__DOT__near_mem$EN_dmem_req = RTL__RTL__DOT__near_mem$EN_dmem_req;
    assign RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL__RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__rg_cur_priv = RTL__RTL__DOT__rg_cur_priv;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    assign RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL__RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL__RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL__RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__DOT__near_mem$dmem_req_addr = RTL__RTL__DOT__near_mem$dmem_req_addr;
    assign RTL__DOT__near_mem$imem_instr = RTL__RTL__DOT__near_mem$imem_instr;
    assign RTL__DOT__f_reset_reqs__DOT__full_reg = RTL__RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__near_mem$imem_pc = RTL__RTL__DOT__near_mem$imem_pc;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem$dmem_exc = RTL__RTL__DOT__near_mem$dmem_exc;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL__RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__DOT__s3_deq$D_IN = RTL__RTL__DOT__s3_deq$D_IN;
    assign RTL__CLK = clk;
    assign RTL__RST_N = ~rst;
    assign RTL__hart0_server_reset_request_put = __VLG_I_hart0_server_reset_request_put;
    assign RTL__EN_hart0_server_reset_request_put = __VLG_I_EN_hart0_server_reset_request_put;
    assign __VLG_O_RDY_hart0_server_reset_request_put = RTL__RDY_hart0_server_reset_request_put;
    assign RTL__EN_hart0_server_reset_response_get = __VLG_I_EN_hart0_server_reset_response_get;
    assign __VLG_O_hart0_server_reset_response_get = RTL__hart0_server_reset_response_get;
    assign __VLG_O_RDY_hart0_server_reset_response_get = RTL__RDY_hart0_server_reset_response_get;
    assign __VLG_O_imem_master_awvalid = RTL__imem_master_awvalid;
    assign __VLG_O_imem_master_awid = RTL__imem_master_awid;
    assign __VLG_O_imem_master_awaddr = RTL__imem_master_awaddr;
    assign __VLG_O_imem_master_awlen = RTL__imem_master_awlen;
    assign __VLG_O_imem_master_awsize = RTL__imem_master_awsize;
    assign __VLG_O_imem_master_awburst = RTL__imem_master_awburst;
    assign __VLG_O_imem_master_awlock = RTL__imem_master_awlock;
    assign __VLG_O_imem_master_awcache = RTL__imem_master_awcache;
    assign __VLG_O_imem_master_awprot = RTL__imem_master_awprot;
    assign __VLG_O_imem_master_awqos = RTL__imem_master_awqos;
    assign __VLG_O_imem_master_awregion = RTL__imem_master_awregion;
    assign RTL__imem_master_awready = __VLG_I_imem_master_awready;
    assign __VLG_O_imem_master_wvalid = RTL__imem_master_wvalid;
    assign __VLG_O_imem_master_wdata = RTL__imem_master_wdata;
    assign __VLG_O_imem_master_wstrb = RTL__imem_master_wstrb;
    assign __VLG_O_imem_master_wlast = RTL__imem_master_wlast;
    assign RTL__imem_master_wready = __VLG_I_imem_master_wready;
    assign RTL__imem_master_bvalid = __VLG_I_imem_master_bvalid;
    assign RTL__imem_master_bid = __VLG_I_imem_master_bid;
    assign RTL__imem_master_bresp = __VLG_I_imem_master_bresp;
    assign __VLG_O_imem_master_bready = RTL__imem_master_bready;
    assign __VLG_O_imem_master_arvalid = RTL__imem_master_arvalid;
    assign __VLG_O_imem_master_arid = RTL__imem_master_arid;
    assign __VLG_O_imem_master_araddr = RTL__imem_master_araddr;
    assign __VLG_O_imem_master_arlen = RTL__imem_master_arlen;
    assign __VLG_O_imem_master_arsize = RTL__imem_master_arsize;
    assign __VLG_O_imem_master_arburst = RTL__imem_master_arburst;
    assign __VLG_O_imem_master_arlock = RTL__imem_master_arlock;
    assign __VLG_O_imem_master_arcache = RTL__imem_master_arcache;
    assign __VLG_O_imem_master_arprot = RTL__imem_master_arprot;
    assign __VLG_O_imem_master_arqos = RTL__imem_master_arqos;
    assign __VLG_O_imem_master_arregion = RTL__imem_master_arregion;
    assign RTL__imem_master_arready = __VLG_I_imem_master_arready;
    assign RTL__imem_master_rvalid = __VLG_I_imem_master_rvalid;
    assign RTL__imem_master_rid = __VLG_I_imem_master_rid;
    assign RTL__imem_master_rdata = __VLG_I_imem_master_rdata;
    assign RTL__imem_master_rresp = __VLG_I_imem_master_rresp;
    assign RTL__imem_master_rlast = __VLG_I_imem_master_rlast;
    assign __VLG_O_imem_master_rready = RTL__imem_master_rready;
    assign __VLG_O_dmem_master_awvalid = RTL__dmem_master_awvalid;
    assign __VLG_O_dmem_master_awid = RTL__dmem_master_awid;
    assign __VLG_O_dmem_master_awaddr = RTL__dmem_master_awaddr;
    assign __VLG_O_dmem_master_awlen = RTL__dmem_master_awlen;
    assign __VLG_O_dmem_master_awsize = RTL__dmem_master_awsize;
    assign __VLG_O_dmem_master_awburst = RTL__dmem_master_awburst;
    assign __VLG_O_dmem_master_awlock = RTL__dmem_master_awlock;
    assign __VLG_O_dmem_master_awcache = RTL__dmem_master_awcache;
    assign __VLG_O_dmem_master_awprot = RTL__dmem_master_awprot;
    assign __VLG_O_dmem_master_awqos = RTL__dmem_master_awqos;
    assign __VLG_O_dmem_master_awregion = RTL__dmem_master_awregion;
    assign RTL__dmem_master_awready = __VLG_I_dmem_master_awready;
    assign __VLG_O_dmem_master_wvalid = RTL__dmem_master_wvalid;
    assign __VLG_O_dmem_master_wdata = RTL__dmem_master_wdata;
    assign __VLG_O_dmem_master_wstrb = RTL__dmem_master_wstrb;
    assign __VLG_O_dmem_master_wlast = RTL__dmem_master_wlast;
    assign RTL__dmem_master_wready = __VLG_I_dmem_master_wready;
    assign RTL__dmem_master_bvalid = __VLG_I_dmem_master_bvalid;
    assign RTL__dmem_master_bid = __VLG_I_dmem_master_bid;
    assign RTL__dmem_master_bresp = __VLG_I_dmem_master_bresp;
    assign __VLG_O_dmem_master_bready = RTL__dmem_master_bready;
    assign __VLG_O_dmem_master_arvalid = RTL__dmem_master_arvalid;
    assign __VLG_O_dmem_master_arid = RTL__dmem_master_arid;
    assign __VLG_O_dmem_master_araddr = RTL__dmem_master_araddr;
    assign __VLG_O_dmem_master_arlen = RTL__dmem_master_arlen;
    assign __VLG_O_dmem_master_arsize = RTL__dmem_master_arsize;
    assign __VLG_O_dmem_master_arburst = RTL__dmem_master_arburst;
    assign __VLG_O_dmem_master_arlock = RTL__dmem_master_arlock;
    assign __VLG_O_dmem_master_arcache = RTL__dmem_master_arcache;
    assign __VLG_O_dmem_master_arprot = RTL__dmem_master_arprot;
    assign __VLG_O_dmem_master_arqos = RTL__dmem_master_arqos;
    assign __VLG_O_dmem_master_arregion = RTL__dmem_master_arregion;
    assign RTL__dmem_master_arready = __VLG_I_dmem_master_arready;
    assign RTL__dmem_master_rvalid = __VLG_I_dmem_master_rvalid;
    assign RTL__dmem_master_rid = __VLG_I_dmem_master_rid;
    assign RTL__dmem_master_rdata = __VLG_I_dmem_master_rdata;
    assign RTL__dmem_master_rresp = __VLG_I_dmem_master_rresp;
    assign RTL__dmem_master_rlast = __VLG_I_dmem_master_rlast;
    assign __VLG_O_dmem_master_rready = RTL__dmem_master_rready;
    assign RTL__m_external_interrupt_req_set_not_clear = __VLG_II_m_external_interrupt_req_set_not_clear;
    assign RTL__s_external_interrupt_req_set_not_clear = __VLG_II_s_external_interrupt_req_set_not_clear;
    assign RTL__software_interrupt_req_set_not_clear = __VLG_II_software_interrupt_req_set_not_clear;
    assign RTL__timer_interrupt_req_set_not_clear = __VLG_II_timer_interrupt_req_set_not_clear;
    assign RTL__nmi_req_set_not_clear = __VLG_II_nmi_req_set_not_clear;
    assign RTL__set_verbosity_verbosity = __VLG_I_set_verbosity_verbosity;
    assign RTL__set_verbosity_logdelay = __VLG_I_set_verbosity_logdelay;
    assign RTL__EN_set_verbosity = __VLG_I_EN_set_verbosity;
    assign __VLG_O_RDY_set_verbosity = RTL__RDY_set_verbosity;
    
assign __all_assert_wire__ = (variable_map_assert__p118__) && (variable_map_assert__p119__) && (variable_map_assert__p120__) && (variable_map_assert__p121__) && (variable_map_assert__p122__) && (variable_map_assert__p123__) && (variable_map_assert__p124__) && (variable_map_assert__p125__) && (variable_map_assert__p126__) && (variable_map_assert__p127__) && (variable_map_assert__p128__) && (variable_map_assert__p129__) && (variable_map_assert__p130__) && (variable_map_assert__p131__) && (variable_map_assert__p132__) && (variable_map_assert__p133__) && (variable_map_assert__p134__) && (variable_map_assert__p135__) && (variable_map_assert__p136__) && (variable_map_assert__p137__) && (variable_map_assert__p138__) && (variable_map_assert__p139__) && (variable_map_assert__p140__) && (variable_map_assert__p141__) && (variable_map_assert__p142__) && (variable_map_assert__p143__) && (variable_map_assert__p144__) && (variable_map_assert__p145__) && (variable_map_assert__p146__) && (variable_map_assert__p147__) && (variable_map_assert__p148__) && (variable_map_assert__p149__) && (variable_map_assert__p150__) && (variable_map_assert__p151__) && (variable_map_assert__p152__) ;
normalassert: assert property ( __all_assert_wire__ ); // the only assertion 

assign __all_assume_wire__ = (input_map_assume___p0__)&& (invariant_assume__p1__)&& (invariant_assume__p2__)&& (invariant_assume__p3__)&& (invariant_assume__p4__)&& (invariant_assume__p5__)&& (invariant_assume__p6__)&& (invariant_assume__p7__)&& (invariant_assume__p8__)&& (invariant_assume__p9__)&& (invariant_assume__p10__)&& (invariant_assume__p11__)&& (invariant_assume__p12__)&& (invariant_assume__p13__)&& (invariant_assume__p14__)&& (invariant_assume__p15__)&& (invariant_assume__p16__)&& (invariant_assume__p17__)&& (invariant_assume__p18__)&& (invariant_assume__p19__)&& (invariant_assume__p20__)&& (invariant_assume__p21__)&& (invariant_assume__p22__)&& (invariant_assume__p23__)&& (invariant_assume__p24__)&& (invariant_assume__p25__)&& (invariant_assume__p26__)&& (invariant_assume__p27__)&& (invariant_assume__p28__)&& (invariant_assume__p29__)&& (invariant_assume__p30__)&& (invariant_assume__p31__)&& (invariant_assume__p32__)&& (issue_decode__p33__)&& (issue_valid__p34__)&& (noreset__p35__)&& (post_value_holder__p36__)&& (post_value_holder__p37__)&& (post_value_holder__p38__)&& (post_value_holder__p39__)&& (post_value_holder__p40__)&& (post_value_holder__p41__)&& (post_value_holder__p42__)&& (post_value_holder__p43__)&& (post_value_holder__p44__)&& (post_value_holder__p45__)&& (post_value_holder__p46__)&& (post_value_holder__p47__)&& (post_value_holder__p48__)&& (post_value_holder__p49__)&& (post_value_holder__p50__)&& (post_value_holder__p51__)&& (post_value_holder__p52__)&& (post_value_holder__p53__)&& (post_value_holder__p54__)&& (post_value_holder__p55__)&& (post_value_holder__p56__)&& (post_value_holder__p57__)&& (post_value_holder__p58__)&& (post_value_holder__p59__)&& (post_value_holder__p60__)&& (post_value_holder__p61__)&& (post_value_holder__p62__)&& (post_value_holder__p63__)&& (post_value_holder__p64__)&& (post_value_holder__p65__)&& (post_value_holder__p66__)&& (post_value_holder__p67__)&& (post_value_holder__p68__)&& (post_value_holder__p69__)&& (post_value_holder__p70__)&& (post_value_holder__p71__)&& (post_value_holder__p72__)&& (post_value_holder__p73__)&& (rfassumptions__p74__)&& (rfassumptions__p75__)&& (rfassumptions__p76__)&& (variable_map_assume___p77__)&& (variable_map_assume___p78__)&& (variable_map_assume___p79__)&& (variable_map_assume___p80__)&& (variable_map_assume___p81__)&& (variable_map_assume___p82__)&& (variable_map_assume___p83__)&& (variable_map_assume___p84__)&& (variable_map_assume___p85__)&& (variable_map_assume___p86__)&& (variable_map_assume___p87__)&& (variable_map_assume___p88__)&& (variable_map_assume___p89__)&& (variable_map_assume___p90__)&& (variable_map_assume___p91__)&& (variable_map_assume___p92__)&& (variable_map_assume___p93__)&& (variable_map_assume___p94__)&& (variable_map_assume___p95__)&& (variable_map_assume___p96__)&& (variable_map_assume___p97__)&& (variable_map_assume___p98__)&& (variable_map_assume___p99__)&& (variable_map_assume___p100__)&& (variable_map_assume___p101__)&& (variable_map_assume___p102__)&& (variable_map_assume___p103__)&& (variable_map_assume___p104__)&& (variable_map_assume___p105__)&& (variable_map_assume___p106__)&& (variable_map_assume___p107__)&& (variable_map_assume___p108__)&& (variable_map_assume___p109__)&& (variable_map_assume___p110__)&& (variable_map_assume___p111__)&& (variable_map_assume___p112__)&& (variable_map_assume___p113__)&& (variable_map_assume___p114__)&& (variable_map_assume___p115__)&& (variable_map_assume___p116__)&& (variable_map_assume___p117__) ;
all_assume: assume property ( __all_assume_wire__ ); // the only sanity assertion 

assign __sanitycheck_wire__ = (post_value_holder_overly_constrained__p153__) && (post_value_holder_overly_constrained__p154__) && (post_value_holder_overly_constrained__p155__) && (post_value_holder_overly_constrained__p156__) && (post_value_holder_overly_constrained__p157__) && (post_value_holder_overly_constrained__p158__) && (post_value_holder_overly_constrained__p159__) && (post_value_holder_overly_constrained__p160__) && (post_value_holder_overly_constrained__p161__) && (post_value_holder_overly_constrained__p162__) && (post_value_holder_overly_constrained__p163__) && (post_value_holder_overly_constrained__p164__) && (post_value_holder_overly_constrained__p165__) && (post_value_holder_overly_constrained__p166__) && (post_value_holder_overly_constrained__p167__) && (post_value_holder_overly_constrained__p168__) && (post_value_holder_overly_constrained__p169__) && (post_value_holder_overly_constrained__p170__) && (post_value_holder_overly_constrained__p171__) && (post_value_holder_overly_constrained__p172__) && (post_value_holder_overly_constrained__p173__) && (post_value_holder_overly_constrained__p174__) && (post_value_holder_overly_constrained__p175__) && (post_value_holder_overly_constrained__p176__) && (post_value_holder_overly_constrained__p177__) && (post_value_holder_overly_constrained__p178__) && (post_value_holder_overly_constrained__p179__) && (post_value_holder_overly_constrained__p180__) && (post_value_holder_overly_constrained__p181__) && (post_value_holder_overly_constrained__p182__) && (post_value_holder_overly_constrained__p183__) && (post_value_holder_overly_constrained__p184__) && (post_value_holder_overly_constrained__p185__) && (post_value_holder_overly_constrained__p186__) && (post_value_holder_overly_constrained__p187__) && (post_value_holder_overly_constrained__p188__) && (post_value_holder_overly_constrained__p189__) && (post_value_holder_overly_constrained__p190__) && (post_value_holder_triggered__p191__) && (post_value_holder_triggered__p192__) && (post_value_holder_triggered__p193__) && (post_value_holder_triggered__p194__) && (post_value_holder_triggered__p195__) && (post_value_holder_triggered__p196__) && (post_value_holder_triggered__p197__) && (post_value_holder_triggered__p198__) && (post_value_holder_triggered__p199__) && (post_value_holder_triggered__p200__) && (post_value_holder_triggered__p201__) && (post_value_holder_triggered__p202__) && (post_value_holder_triggered__p203__) && (post_value_holder_triggered__p204__) && (post_value_holder_triggered__p205__) && (post_value_holder_triggered__p206__) && (post_value_holder_triggered__p207__) && (post_value_holder_triggered__p208__) && (post_value_holder_triggered__p209__) && (post_value_holder_triggered__p210__) && (post_value_holder_triggered__p211__) && (post_value_holder_triggered__p212__) && (post_value_holder_triggered__p213__) && (post_value_holder_triggered__p214__) && (post_value_holder_triggered__p215__) && (post_value_holder_triggered__p216__) && (post_value_holder_triggered__p217__) && (post_value_holder_triggered__p218__) && (post_value_holder_triggered__p219__) && (post_value_holder_triggered__p220__) && (post_value_holder_triggered__p221__) && (post_value_holder_triggered__p222__) && (post_value_holder_triggered__p223__) && (post_value_holder_triggered__p224__) && (post_value_holder_triggered__p225__) && (post_value_holder_triggered__p226__) && (post_value_holder_triggered__p227__) && (post_value_holder_triggered__p228__) ;
sanitycheck: assert property ( __sanitycheck_wire__ ); // the only assumption 

always @(posedge clk) begin
   if(rst) begin
       __auxvar10__recorder <= ____auxvar10__recorder_init__;
       __auxvar10__recorder_sn_condmet <= 1'b0;
       __auxvar11__recorder <= ____auxvar11__recorder_init__;
       __auxvar11__recorder_sn_condmet <= 1'b0;
       __auxvar12__recorder <= ____auxvar12__recorder_init__;
       __auxvar12__recorder_sn_condmet <= 1'b0;
       __auxvar13__recorder <= ____auxvar13__recorder_init__;
       __auxvar13__recorder_sn_condmet <= 1'b0;
       __auxvar14__recorder <= ____auxvar14__recorder_init__;
       __auxvar14__recorder_sn_condmet <= 1'b0;
       __auxvar15__recorder <= ____auxvar15__recorder_init__;
       __auxvar15__recorder_sn_condmet <= 1'b0;
       __auxvar16__recorder <= ____auxvar16__recorder_init__;
       __auxvar16__recorder_sn_condmet <= 1'b0;
       __auxvar17__recorder <= ____auxvar17__recorder_init__;
       __auxvar17__recorder_sn_condmet <= 1'b0;
       __auxvar18__recorder <= ____auxvar18__recorder_init__;
       __auxvar18__recorder_sn_condmet <= 1'b0;
       __auxvar19__recorder <= ____auxvar19__recorder_init__;
       __auxvar19__recorder_sn_condmet <= 1'b0;
       __auxvar1__recorder <= ____auxvar1__recorder_init__;
       __auxvar1__recorder_sn_condmet <= 1'b0;
       __auxvar20__recorder <= ____auxvar20__recorder_init__;
       __auxvar20__recorder_sn_condmet <= 1'b0;
       __auxvar21__recorder <= ____auxvar21__recorder_init__;
       __auxvar21__recorder_sn_condmet <= 1'b0;
       __auxvar22__recorder <= ____auxvar22__recorder_init__;
       __auxvar22__recorder_sn_condmet <= 1'b0;
       __auxvar23__recorder <= ____auxvar23__recorder_init__;
       __auxvar23__recorder_sn_condmet <= 1'b0;
       __auxvar24__recorder <= ____auxvar24__recorder_init__;
       __auxvar24__recorder_sn_condmet <= 1'b0;
       __auxvar25__recorder <= ____auxvar25__recorder_init__;
       __auxvar25__recorder_sn_condmet <= 1'b0;
       __auxvar26__recorder <= ____auxvar26__recorder_init__;
       __auxvar26__recorder_sn_condmet <= 1'b0;
       __auxvar27__recorder <= ____auxvar27__recorder_init__;
       __auxvar27__recorder_sn_condmet <= 1'b0;
       __auxvar28__recorder <= ____auxvar28__recorder_init__;
       __auxvar28__recorder_sn_condmet <= 1'b0;
       __auxvar29__recorder <= ____auxvar29__recorder_init__;
       __auxvar29__recorder_sn_condmet <= 1'b0;
       __auxvar2__recorder <= ____auxvar2__recorder_init__;
       __auxvar2__recorder_sn_condmet <= 1'b0;
       __auxvar30__recorder <= ____auxvar30__recorder_init__;
       __auxvar30__recorder_sn_condmet <= 1'b0;
       __auxvar31__recorder <= ____auxvar31__recorder_init__;
       __auxvar31__recorder_sn_condmet <= 1'b0;
       __auxvar32__recorder <= ____auxvar32__recorder_init__;
       __auxvar32__recorder_sn_condmet <= 1'b0;
       __auxvar33__recorder <= ____auxvar33__recorder_init__;
       __auxvar33__recorder_sn_condmet <= 1'b0;
       __auxvar34__recorder <= ____auxvar34__recorder_init__;
       __auxvar34__recorder_sn_condmet <= 1'b0;
       __auxvar35__recorder <= ____auxvar35__recorder_init__;
       __auxvar35__recorder_sn_condmet <= 1'b0;
       __auxvar36__recorder <= ____auxvar36__recorder_init__;
       __auxvar36__recorder_sn_condmet <= 1'b0;
       __auxvar37__recorder <= ____auxvar37__recorder_init__;
       __auxvar37__recorder_sn_condmet <= 1'b0;
       __auxvar38__recorder <= ____auxvar38__recorder_init__;
       __auxvar38__recorder_sn_condmet <= 1'b0;
       __auxvar3__recorder <= ____auxvar3__recorder_init__;
       __auxvar3__recorder_sn_condmet <= 1'b0;
       __auxvar4__recorder <= ____auxvar4__recorder_init__;
       __auxvar4__recorder_sn_condmet <= 1'b0;
       __auxvar5__recorder <= ____auxvar5__recorder_init__;
       __auxvar5__recorder_sn_condmet <= 1'b0;
       __auxvar6__recorder <= ____auxvar6__recorder_init__;
       __auxvar6__recorder_sn_condmet <= 1'b0;
       __auxvar7__recorder <= ____auxvar7__recorder_init__;
       __auxvar7__recorder_sn_condmet <= 1'b0;
       __auxvar8__recorder <= ____auxvar8__recorder_init__;
       __auxvar8__recorder_sn_condmet <= 1'b0;
       __auxvar9__recorder <= ____auxvar9__recorder_init__;
       __auxvar9__recorder_sn_condmet <= 1'b0;
       __auxvar0__delay_d_1<= 0;
       monitor_s1_already<= 1'b0;
       monitor_s2<= 1'b0;
       monitor_s3<= 1'b0;
       monitor_s4<= 1'b0;
   end
   else if(1) begin
       __auxvar10__recorder <= __auxvar10__recorder;
       if (__auxvar10__recorder_sn_cond ) begin __auxvar10__recorder_sn_condmet <= 1'b1; __auxvar10__recorder_sn_vhold <= __auxvar10__recorder_sn_value; end
       __auxvar11__recorder <= __auxvar11__recorder;
       if (__auxvar11__recorder_sn_cond ) begin __auxvar11__recorder_sn_condmet <= 1'b1; __auxvar11__recorder_sn_vhold <= __auxvar11__recorder_sn_value; end
       __auxvar12__recorder <= __auxvar12__recorder;
       if (__auxvar12__recorder_sn_cond ) begin __auxvar12__recorder_sn_condmet <= 1'b1; __auxvar12__recorder_sn_vhold <= __auxvar12__recorder_sn_value; end
       __auxvar13__recorder <= __auxvar13__recorder;
       if (__auxvar13__recorder_sn_cond ) begin __auxvar13__recorder_sn_condmet <= 1'b1; __auxvar13__recorder_sn_vhold <= __auxvar13__recorder_sn_value; end
       __auxvar14__recorder <= __auxvar14__recorder;
       if (__auxvar14__recorder_sn_cond ) begin __auxvar14__recorder_sn_condmet <= 1'b1; __auxvar14__recorder_sn_vhold <= __auxvar14__recorder_sn_value; end
       __auxvar15__recorder <= __auxvar15__recorder;
       if (__auxvar15__recorder_sn_cond ) begin __auxvar15__recorder_sn_condmet <= 1'b1; __auxvar15__recorder_sn_vhold <= __auxvar15__recorder_sn_value; end
       __auxvar16__recorder <= __auxvar16__recorder;
       if (__auxvar16__recorder_sn_cond ) begin __auxvar16__recorder_sn_condmet <= 1'b1; __auxvar16__recorder_sn_vhold <= __auxvar16__recorder_sn_value; end
       __auxvar17__recorder <= __auxvar17__recorder;
       if (__auxvar17__recorder_sn_cond ) begin __auxvar17__recorder_sn_condmet <= 1'b1; __auxvar17__recorder_sn_vhold <= __auxvar17__recorder_sn_value; end
       __auxvar18__recorder <= __auxvar18__recorder;
       if (__auxvar18__recorder_sn_cond ) begin __auxvar18__recorder_sn_condmet <= 1'b1; __auxvar18__recorder_sn_vhold <= __auxvar18__recorder_sn_value; end
       __auxvar19__recorder <= __auxvar19__recorder;
       if (__auxvar19__recorder_sn_cond ) begin __auxvar19__recorder_sn_condmet <= 1'b1; __auxvar19__recorder_sn_vhold <= __auxvar19__recorder_sn_value; end
       __auxvar1__recorder <= __auxvar1__recorder;
       if (__auxvar1__recorder_sn_cond ) begin __auxvar1__recorder_sn_condmet <= 1'b1; __auxvar1__recorder_sn_vhold <= __auxvar1__recorder_sn_value; end
       __auxvar20__recorder <= __auxvar20__recorder;
       if (__auxvar20__recorder_sn_cond ) begin __auxvar20__recorder_sn_condmet <= 1'b1; __auxvar20__recorder_sn_vhold <= __auxvar20__recorder_sn_value; end
       __auxvar21__recorder <= __auxvar21__recorder;
       if (__auxvar21__recorder_sn_cond ) begin __auxvar21__recorder_sn_condmet <= 1'b1; __auxvar21__recorder_sn_vhold <= __auxvar21__recorder_sn_value; end
       __auxvar22__recorder <= __auxvar22__recorder;
       if (__auxvar22__recorder_sn_cond ) begin __auxvar22__recorder_sn_condmet <= 1'b1; __auxvar22__recorder_sn_vhold <= __auxvar22__recorder_sn_value; end
       __auxvar23__recorder <= __auxvar23__recorder;
       if (__auxvar23__recorder_sn_cond ) begin __auxvar23__recorder_sn_condmet <= 1'b1; __auxvar23__recorder_sn_vhold <= __auxvar23__recorder_sn_value; end
       __auxvar24__recorder <= __auxvar24__recorder;
       if (__auxvar24__recorder_sn_cond ) begin __auxvar24__recorder_sn_condmet <= 1'b1; __auxvar24__recorder_sn_vhold <= __auxvar24__recorder_sn_value; end
       __auxvar25__recorder <= __auxvar25__recorder;
       if (__auxvar25__recorder_sn_cond ) begin __auxvar25__recorder_sn_condmet <= 1'b1; __auxvar25__recorder_sn_vhold <= __auxvar25__recorder_sn_value; end
       __auxvar26__recorder <= __auxvar26__recorder;
       if (__auxvar26__recorder_sn_cond ) begin __auxvar26__recorder_sn_condmet <= 1'b1; __auxvar26__recorder_sn_vhold <= __auxvar26__recorder_sn_value; end
       __auxvar27__recorder <= __auxvar27__recorder;
       if (__auxvar27__recorder_sn_cond ) begin __auxvar27__recorder_sn_condmet <= 1'b1; __auxvar27__recorder_sn_vhold <= __auxvar27__recorder_sn_value; end
       __auxvar28__recorder <= __auxvar28__recorder;
       if (__auxvar28__recorder_sn_cond ) begin __auxvar28__recorder_sn_condmet <= 1'b1; __auxvar28__recorder_sn_vhold <= __auxvar28__recorder_sn_value; end
       __auxvar29__recorder <= __auxvar29__recorder;
       if (__auxvar29__recorder_sn_cond ) begin __auxvar29__recorder_sn_condmet <= 1'b1; __auxvar29__recorder_sn_vhold <= __auxvar29__recorder_sn_value; end
       __auxvar2__recorder <= __auxvar2__recorder;
       if (__auxvar2__recorder_sn_cond ) begin __auxvar2__recorder_sn_condmet <= 1'b1; __auxvar2__recorder_sn_vhold <= __auxvar2__recorder_sn_value; end
       __auxvar30__recorder <= __auxvar30__recorder;
       if (__auxvar30__recorder_sn_cond ) begin __auxvar30__recorder_sn_condmet <= 1'b1; __auxvar30__recorder_sn_vhold <= __auxvar30__recorder_sn_value; end
       __auxvar31__recorder <= __auxvar31__recorder;
       if (__auxvar31__recorder_sn_cond ) begin __auxvar31__recorder_sn_condmet <= 1'b1; __auxvar31__recorder_sn_vhold <= __auxvar31__recorder_sn_value; end
       __auxvar32__recorder <= __auxvar32__recorder;
       if (__auxvar32__recorder_sn_cond ) begin __auxvar32__recorder_sn_condmet <= 1'b1; __auxvar32__recorder_sn_vhold <= __auxvar32__recorder_sn_value; end
       __auxvar33__recorder <= __auxvar33__recorder;
       if (__auxvar33__recorder_sn_cond ) begin __auxvar33__recorder_sn_condmet <= 1'b1; __auxvar33__recorder_sn_vhold <= __auxvar33__recorder_sn_value; end
       __auxvar34__recorder <= __auxvar34__recorder;
       if (__auxvar34__recorder_sn_cond ) begin __auxvar34__recorder_sn_condmet <= 1'b1; __auxvar34__recorder_sn_vhold <= __auxvar34__recorder_sn_value; end
       __auxvar35__recorder <= __auxvar35__recorder;
       if (__auxvar35__recorder_sn_cond ) begin __auxvar35__recorder_sn_condmet <= 1'b1; __auxvar35__recorder_sn_vhold <= __auxvar35__recorder_sn_value; end
       __auxvar36__recorder <= __auxvar36__recorder;
       if (__auxvar36__recorder_sn_cond ) begin __auxvar36__recorder_sn_condmet <= 1'b1; __auxvar36__recorder_sn_vhold <= __auxvar36__recorder_sn_value; end
       __auxvar37__recorder <= __auxvar37__recorder;
       if (__auxvar37__recorder_sn_cond ) begin __auxvar37__recorder_sn_condmet <= 1'b1; __auxvar37__recorder_sn_vhold <= __auxvar37__recorder_sn_value; end
       __auxvar38__recorder <= __auxvar38__recorder;
       if (__auxvar38__recorder_sn_cond ) begin __auxvar38__recorder_sn_condmet <= 1'b1; __auxvar38__recorder_sn_vhold <= __auxvar38__recorder_sn_value; end
       __auxvar3__recorder <= __auxvar3__recorder;
       if (__auxvar3__recorder_sn_cond ) begin __auxvar3__recorder_sn_condmet <= 1'b1; __auxvar3__recorder_sn_vhold <= __auxvar3__recorder_sn_value; end
       __auxvar4__recorder <= __auxvar4__recorder;
       if (__auxvar4__recorder_sn_cond ) begin __auxvar4__recorder_sn_condmet <= 1'b1; __auxvar4__recorder_sn_vhold <= __auxvar4__recorder_sn_value; end
       __auxvar5__recorder <= __auxvar5__recorder;
       if (__auxvar5__recorder_sn_cond ) begin __auxvar5__recorder_sn_condmet <= 1'b1; __auxvar5__recorder_sn_vhold <= __auxvar5__recorder_sn_value; end
       __auxvar6__recorder <= __auxvar6__recorder;
       if (__auxvar6__recorder_sn_cond ) begin __auxvar6__recorder_sn_condmet <= 1'b1; __auxvar6__recorder_sn_vhold <= __auxvar6__recorder_sn_value; end
       __auxvar7__recorder <= __auxvar7__recorder;
       if (__auxvar7__recorder_sn_cond ) begin __auxvar7__recorder_sn_condmet <= 1'b1; __auxvar7__recorder_sn_vhold <= __auxvar7__recorder_sn_value; end
       __auxvar8__recorder <= __auxvar8__recorder;
       if (__auxvar8__recorder_sn_cond ) begin __auxvar8__recorder_sn_condmet <= 1'b1; __auxvar8__recorder_sn_vhold <= __auxvar8__recorder_sn_value; end
       __auxvar9__recorder <= __auxvar9__recorder;
       if (__auxvar9__recorder_sn_cond ) begin __auxvar9__recorder_sn_condmet <= 1'b1; __auxvar9__recorder_sn_vhold <= __auxvar9__recorder_sn_value; end
       __auxvar0__delay_d_1 <= __auxvar0__delay_d_0 ;
       if(monitor_s1_already_enter_cond) begin monitor_s1_already <= 1'b1;
       end
       else if(monitor_s1_already_exit_cond) begin monitor_s1_already <= 1'b0;
       end
       if(monitor_s2_enter_cond) begin monitor_s2 <= 1'b1;
       end
       else if(monitor_s2_exit_cond) begin monitor_s2 <= 1'b0;
       end
       if(monitor_s3_enter_cond) begin monitor_s3 <= 1'b1;
       end
       else if(monitor_s3_exit_cond) begin monitor_s3 <= 1'b0;
       end
       if(monitor_s4_enter_cond) begin monitor_s4 <= 1'b1;
       end
       else if(monitor_s4_exit_cond) begin monitor_s4 <= 1'b0;
       end
   end
end
endmodule