module RocketTile(
  input         clock,
                reset,
  output        auto_buffer_in_a_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_in_a_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [2:0]  auto_buffer_in_a_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_in_a_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_in_a_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [4:0]  auto_buffer_in_a_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [31:0] auto_buffer_in_a_bits_address,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [3:0]  auto_buffer_in_a_bits_mask,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [31:0] auto_buffer_in_a_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_in_a_bits_corrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_in_d_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_in_d_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [2:0]  auto_buffer_in_d_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_in_d_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [4:0]  auto_buffer_in_d_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_buffer_in_d_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_a_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_a_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [2:0]  auto_buffer_out_a_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [3:0]  auto_buffer_out_a_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_a_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_buffer_out_a_bits_address,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [3:0]  auto_buffer_out_a_bits_mask,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_buffer_out_a_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_d_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_d_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [2:0]  auto_buffer_out_d_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [1:0]  auto_buffer_out_d_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [3:0]  auto_buffer_out_d_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_d_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_d_bits_sink,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_d_bits_denied,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [31:0] auto_buffer_out_d_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_d_bits_corrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_broadcast_out_insns_0_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_broadcast_out_insns_0_iaddr,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_broadcast_out_insns_0_insn,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [2:0]  auto_broadcast_out_insns_0_priv,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_broadcast_out_insns_0_exception,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_broadcast_out_insns_0_interrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_broadcast_out_insns_0_cause,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_broadcast_out_insns_0_tval,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [63:0] auto_broadcast_out_time,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_wfi_out_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_int_local_in_2_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_int_local_in_1_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_int_local_in_1_1,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_int_local_in_0_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_hartid_in	// src/main/scala/diplomacy/LazyModule.scala:374:18
);

  wire        intSinkNodeIn_3;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        intSinkNodeIn_2;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        intSinkNodeIn_1;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        intSinkNodeIn_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] buffer_1_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [4:0]  buffer_1_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_1_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_1_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_1_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_1_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_1_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_1_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_1_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_1_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [4:0]  buffer_1_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_1_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_1_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_1_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_1_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_1_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] widget_1_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_1_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_1_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_1_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] widget_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_nodeIn_time;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] broadcast_3_nodeIn_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] broadcast_3_nodeIn_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_3_nodeIn_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_3_nodeIn_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  broadcast_3_nodeIn_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] broadcast_3_nodeIn_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] broadcast_3_nodeIn_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_3_nodeIn_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlSlaveXbar_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [4:0]  tlSlaveXbar_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  tlSlaveXbar_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  tlSlaveXbar_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlSlaveXbar_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlSlaveXbar_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] tlSlaveXbar_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [4:0]  tlSlaveXbar_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlSlaveXbar_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlSlaveXbar_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlSlaveXbar_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlSlaveXbar_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlSlaveXbar_nodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlSlaveXbar_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlSlaveXbar_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlSlaveXbar_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [4:0]  tlSlaveXbar_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlSlaveXbar_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlSlaveXbar_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlSlaveXbar_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlSlaveXbar_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlSlaveXbar_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        _core_io_imem_might_request;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_req_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_imem_req_bits_pc;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_req_bits_speculative;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_resp_ready;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_bht_update_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_flush_icache;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_progress;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_dmem_req_bits_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [6:0]  _core_io_dmem_req_bits_tag;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [4:0]  _core_io_dmem_req_bits_cmd;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_dmem_req_bits_size;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_signed;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_dv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_s1_kill;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_dmem_s1_data_data;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_bits_rs1;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_debug;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_0_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_0_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_0_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_1_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_1_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_1_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_2_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_2_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_2_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_3_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_3_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_3_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_4_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_4_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_4_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_5_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_5_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_5_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_6_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_6_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_6_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_7_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_7_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_7_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_customCSRs_csrs_0_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_wfi;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _ptw_io_requestor_0_resp_bits_ae_ptw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_ae_final;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_gf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_hr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_hw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_hx;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_0_resp_bits_pte_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_d;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_g;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_u;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_gpa_is_pte;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_debug;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_0_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_0_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_0_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_1_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_1_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_1_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_2_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_2_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_2_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_3_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_3_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_3_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_4_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_4_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_4_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_5_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_5_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_5_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_6_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_6_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_6_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_7_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_7_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_7_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_ae_ptw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_ae_final;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_gf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_hr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_hw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_hx;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_1_resp_bits_pte_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_d;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_g;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_u;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_gpa_is_pte;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_debug;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_0_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_0_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_0_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_1_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_1_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_1_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_2_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_2_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_2_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_3_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_3_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_3_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_4_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_4_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_4_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_5_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_5_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_5_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_6_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_6_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_6_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_7_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_7_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_7_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_customCSRs_csrs_0_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _dcacheArb_io_requestor_0_req_ready;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_nack;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_valid;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [6:0]  _dcacheArb_io_requestor_0_resp_bits_tag;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [31:0] _dcacheArb_io_requestor_0_resp_bits_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_bits_replay;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_bits_has_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [31:0] _dcacheArb_io_requestor_0_resp_bits_data_word_bypass;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_replay_next;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ma_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ma_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_pf_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_pf_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ae_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ae_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_ordered;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_grant;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_1_req_ready;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_1_s2_nack;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_1_resp_valid;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [31:0] _dcacheArb_io_requestor_1_resp_bits_data_raw;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_valid;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [31:0] _dcacheArb_io_mem_req_bits_addr;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [6:0]  _dcacheArb_io_mem_req_bits_tag;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [4:0]  _dcacheArb_io_mem_req_bits_cmd;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [1:0]  _dcacheArb_io_mem_req_bits_size;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_signed;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [1:0]  _dcacheArb_io_mem_req_bits_dprv;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_dv;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_phys;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_no_xcpt;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_s1_kill;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [31:0] _dcacheArb_io_mem_s1_data_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [3:0]  _dcacheArb_io_mem_s1_data_mask;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _fragmenter_1_auto_out_a_valid;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [2:0]  _fragmenter_1_auto_out_a_bits_opcode;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [2:0]  _fragmenter_1_auto_out_a_bits_param;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [1:0]  _fragmenter_1_auto_out_a_bits_size;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [10:0] _fragmenter_1_auto_out_a_bits_source;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [31:0] _fragmenter_1_auto_out_a_bits_address;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [3:0]  _fragmenter_1_auto_out_a_bits_mask;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire [31:0] _fragmenter_1_auto_out_a_bits_data;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire        _fragmenter_1_auto_out_a_bits_corrupt;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire        _fragmenter_1_auto_out_d_ready;	// src/main/scala/tilelink/Fragmenter.scala:335:34
  wire        _dtim_adapter_auto_in_a_ready;	// src/main/scala/tile/RocketTile.scala:60:15
  wire        _dtim_adapter_auto_in_d_valid;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [2:0]  _dtim_adapter_auto_in_d_bits_opcode;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [1:0]  _dtim_adapter_auto_in_d_bits_size;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [10:0] _dtim_adapter_auto_in_d_bits_source;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [31:0] _dtim_adapter_auto_in_d_bits_data;	// src/main/scala/tile/RocketTile.scala:60:15
  wire        _dtim_adapter_io_dmem_req_valid;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [31:0] _dtim_adapter_io_dmem_req_bits_addr;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [4:0]  _dtim_adapter_io_dmem_req_bits_cmd;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [1:0]  _dtim_adapter_io_dmem_req_bits_size;	// src/main/scala/tile/RocketTile.scala:60:15
  wire        _dtim_adapter_io_dmem_s1_kill;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [31:0] _dtim_adapter_io_dmem_s1_data_data;	// src/main/scala/tile/RocketTile.scala:60:15
  wire [3:0]  _dtim_adapter_io_dmem_s1_data_mask;	// src/main/scala/tile/RocketTile.scala:60:15
  wire        _frontend_io_cpu_resp_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [1:0]  _frontend_io_cpu_resp_bits_btb_cfiType;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_taken;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [1:0]  _frontend_io_cpu_resp_bits_btb_mask;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_bridx;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] _frontend_io_cpu_resp_bits_btb_target;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_entry;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [7:0]  _frontend_io_cpu_resp_bits_btb_bht_history;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_bht_value;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] _frontend_io_cpu_resp_bits_pc;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] _frontend_io_cpu_resp_bits_data;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [1:0]  _frontend_io_cpu_resp_bits_mask;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_xcpt_pf_inst;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_xcpt_gf_inst;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_xcpt_ae_inst;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_replay;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_gpa_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] _frontend_io_cpu_gpa_bits;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [19:0] _frontend_io_ptw_req_bits_bits_addr;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_bits_need_gpa;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_bits_vstage1;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_bits_stage2;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _dcache_io_cpu_req_ready;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_nack;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_valid;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [6:0]  _dcache_io_cpu_resp_bits_tag;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [31:0] _dcache_io_cpu_resp_bits_data;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_bits_replay;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_bits_has_data;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [31:0] _dcache_io_cpu_resp_bits_data_word_bypass;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [31:0] _dcache_io_cpu_resp_bits_data_raw;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_replay_next;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ma_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ma_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_pf_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_pf_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ae_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ae_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_ordered;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_grant;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [19:0] _dcache_io_ptw_req_bits_bits_addr;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_bits_need_gpa;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_bits_vstage1;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_bits_stage2;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        buffer_nodeOut_a_ready = auto_buffer_out_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_valid = auto_buffer_out_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_d_bits_opcode = auto_buffer_out_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_d_bits_param = auto_buffer_out_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_d_bits_size = auto_buffer_out_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_bits_source = auto_buffer_out_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_bits_sink = auto_buffer_out_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_bits_denied = auto_buffer_out_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeOut_d_bits_data = auto_buffer_out_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_bits_corrupt = auto_buffer_out_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_1_nodeIn_a_valid = auto_buffer_in_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_1_nodeIn_a_bits_opcode = auto_buffer_in_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_1_nodeIn_a_bits_param = auto_buffer_in_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_1_nodeIn_a_bits_size = auto_buffer_in_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [4:0]  buffer_1_nodeIn_a_bits_source = auto_buffer_in_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] buffer_1_nodeIn_a_bits_address = auto_buffer_in_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  buffer_1_nodeIn_a_bits_mask = auto_buffer_in_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] buffer_1_nodeIn_a_bits_data = auto_buffer_in_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_1_nodeIn_a_bits_corrupt = auto_buffer_in_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_1_nodeIn_d_ready = auto_buffer_in_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        hartidIn = auto_hartid_in;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        int_localIn_0 = auto_int_local_in_0_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        x1_int_localIn_0 = auto_int_local_in_1_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        x1_int_localIn_1 = auto_int_local_in_1_1;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        x1_int_localIn_1_0 = auto_int_local_in_2_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_1_nodeOut_a_bits_mask = 4'hF;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42
  wire [3:0]  widget_1_nodeIn_a_bits_mask = 4'hF;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42
  wire [1:0]  tlSlaveXbar_nodeOut_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  tlSlaveXbar_nodeIn_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  tlSlaveXbar_in_0_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  tlSlaveXbar_out_0_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  tlSlaveXbar_portsBIO_filtered_0_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  tlSlaveXbar_portsDIO_filtered_0_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  buffer_1_nodeOut_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  buffer_1_nodeIn_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  slaveNodeOut_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [1:0]  slaveNodeIn_d_bits_param = 2'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire [3:0]  tlSlaveXbar_beatsBO_decode = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Edges.scala:221:59
  wire [3:0]  tlSlaveXbar_beatsBO_0 = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Edges.scala:222:14
  wire [3:0]  tlSlaveXbar_beatsCI_decode = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Edges.scala:221:59
  wire [3:0]  tlSlaveXbar_beatsCI_0 = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Edges.scala:222:14
  wire [3:0]  tlSlaveXbar_portsBIO_filtered_0_bits_mask = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Xbar.scala:348:24
  wire [3:0]  traceCoreSourceNodeOut_group_0_itype = 4'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [3:0]  traceCoreSourceNodeOut_priv = 4'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [4:0]  tlSlaveXbar_requestBOI_uncommonBits = 5'h0;	// src/main/scala/diplomacy/Parameters.scala:52:56, src/main/scala/tilelink/Bundles.scala:259:74
  wire [4:0]  tlSlaveXbar_portsBIO_filtered_0_bits_source = 5'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Xbar.scala:348:24
  wire [4:0]  tlSlaveXbar_portsCOI_filtered_0_bits_source = 5'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  widget_1_nodeOut_a_bits_opcode = 3'h4;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42
  wire [2:0]  widget_1_nodeIn_a_bits_opcode = 3'h4;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42
  wire [2:0]  tlSlaveXbar_portsBIO_filtered_0_bits_opcode = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  tlSlaveXbar_portsBIO_filtered_0_bits_size = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  tlSlaveXbar_portsCOI_filtered_0_bits_opcode = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  tlSlaveXbar_portsCOI_filtered_0_bits_param = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  tlSlaveXbar_portsCOI_filtered_0_bits_size = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  widget_1_nodeOut_a_bits_param = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [2:0]  widget_1_nodeIn_a_bits_param = 3'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tilelink/Xbar.scala:348:24
  wire [3:0]  widget_1_nodeOut_a_bits_size = 4'h6;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42
  wire [3:0]  widget_1_nodeIn_a_bits_size = 4'h6;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/tile/BaseTile.scala:218:42
  wire [31:0] broadcast_1_nodeIn = 32'h10040;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] broadcast_1_nodeOut = 32'h10040;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] broadcast_1_x1_nodeOut = 32'h10040;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] resetVectorSinkNodeIn = 32'h10040;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] reset_vectorOut = 32'h10040;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] reset_vectorIn = 32'h10040;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] tlSlaveXbar_portsBIO_filtered_0_bits_address = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] tlSlaveXbar_portsBIO_filtered_0_bits_data = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] tlSlaveXbar_portsCOI_filtered_0_bits_address = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] tlSlaveXbar_portsCOI_filtered_0_bits_data = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] broadcast_2_nodeIn_rnmi_interrupt_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] broadcast_2_nodeIn_rnmi_exception_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] broadcast_2_nodeOut_rnmi_interrupt_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] broadcast_2_nodeOut_rnmi_exception_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] widget_1_nodeOut_a_bits_data = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] widget_1_nodeIn_a_bits_data = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] nmiSinkNodeIn_rnmi_interrupt_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] nmiSinkNodeIn_rnmi_exception_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] nmiOut_rnmi_interrupt_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] nmiOut_rnmi_exception_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] nmiIn_rnmi_interrupt_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] nmiIn_rnmi_exception_vector = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] traceCoreSourceNodeOut_group_0_iaddr = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] traceCoreSourceNodeOut_tval = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire [31:0] traceCoreSourceNodeOut_cause = 32'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Xbar.scala:348:24
  wire        tlSlaveXbar_nodeOut_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_nodeOut_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_nodeOut_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_nodeIn_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_nodeIn_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_nodeIn_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_in_0_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_in_0_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_in_0_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_out_0_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_out_0_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_out_0_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_beatsCI_opdata = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsBIO_filtered_0_ready = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsBIO_filtered_0_valid = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsBIO_filtered_0_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsCOI_filtered_0_ready = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsCOI_filtered_0_valid = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsCOI_filtered_0_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsDIO_filtered_0_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsDIO_filtered_0_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsDIO_filtered_0_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsEOI_filtered_0_ready = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsEOI_filtered_0_valid = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_portsEOI_filtered_0_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        broadcast_2_nodeIn_rnmi = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        broadcast_2_nodeOut_rnmi = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_nodeOut = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_1_x1_bundleOut_x_sourceOpt_enable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_1_x1_bundleOut_x_sourceOpt_stall = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_1_nodeOut_enable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_1_nodeOut_stall = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_1_defaultWireOpt_enable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nexus_1_defaultWireOpt_stall = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        broadcast_4_nodeIn_0_rvalid_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        broadcast_4_nodeIn_0_wvalid_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        broadcast_4_nodeIn_0_ivalid_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeOut_a_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeOut_a_bits_user_amba_prot_fetch = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeOut_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeOut_d_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeIn_a_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeIn_a_bits_user_amba_prot_fetch = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeIn_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_nodeIn_d_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_1_nodeOut_a_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_1_nodeOut_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_1_nodeOut_d_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_1_nodeIn_a_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_1_nodeIn_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        widget_1_nodeIn_d_bits_source = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_bufferable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_modifiable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_readalloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_writealloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_privileged = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_secure = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_user_amba_prot_fetch = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeOut_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_bufferable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_modifiable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_readalloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_writealloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_privileged = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_secure = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_user_amba_prot_fetch = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_nodeIn_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_1_nodeOut_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_1_nodeOut_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_1_nodeOut_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_1_nodeIn_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_1_nodeIn_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        buffer_1_nodeIn_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_bufferable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_modifiable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_readalloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_writealloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_privileged = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_secure = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_fetch = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeOut_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_bufferable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_modifiable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_readalloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_writealloc = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_privileged = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_secure = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_fetch = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlOtherMastersNodeIn_a_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nmiSinkNodeIn_rnmi = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nmiOut_rnmi = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        nmiIn_rnmi = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        traceCoreSourceNodeOut_group_0_iretire = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        traceCoreSourceNodeOut_group_0_ilastsize = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        bundleIn_x_sourceOpt_enable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        bundleIn_x_sourceOpt_stall = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        traceAuxSinkNodeIn_enable = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        traceAuxSinkNodeIn_stall = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        bpwatchSourceNodeOut_0_rvalid_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        bpwatchSourceNodeOut_0_wvalid_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        bpwatchSourceNodeOut_0_ivalid_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        haltNodeOut_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        ceaseNodeOut_0 = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        slaveNodeOut_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        slaveNodeOut_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        slaveNodeOut_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        slaveNodeIn_d_bits_sink = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        slaveNodeIn_d_bits_denied = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        slaveNodeIn_d_bits_corrupt = 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
  wire        tlSlaveXbar_requestAIO_0_0 = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        tlSlaveXbar_requestCIO_0_0 = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        tlSlaveXbar_requestBOI_0_0 = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        tlSlaveXbar_requestDOI_0_0 = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        tlSlaveXbar_beatsBO_opdata = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_nodeOut_a_bits_user_amba_prot_secure = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_nodeIn_a_bits_user_amba_prot_secure = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeOut_a_bits_user_amba_prot_bufferable = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeOut_a_bits_user_amba_prot_modifiable = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeOut_a_bits_user_amba_prot_privileged = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeOut_a_bits_user_amba_prot_secure = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeOut_a_bits_user_amba_prot_fetch = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeOut_d_ready = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeIn_a_bits_user_amba_prot_bufferable = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeIn_a_bits_user_amba_prot_modifiable = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeIn_a_bits_user_amba_prot_privileged = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeIn_a_bits_user_amba_prot_secure = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeIn_a_bits_user_amba_prot_fetch = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        widget_1_nodeIn_d_ready = 1'h1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/diplomacy/Parameters.scala:56:48, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/tile/BaseTile.scala:218:42, src/main/scala/tile/RocketTile.scala:127:20, src/main/scala/tilelink/Edges.scala:98:28, src/main/scala/tilelink/Xbar.scala:303:107, :304:107
  wire        tlSlaveXbar_out_0_a_ready = tlSlaveXbar_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_out_0_a_valid;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_out_0_a_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_out_0_a_bits_param;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_out_0_a_bits_size;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [4:0]  tlSlaveXbar_out_0_a_bits_source;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [31:0] tlSlaveXbar_out_0_a_bits_address;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [3:0]  tlSlaveXbar_out_0_a_bits_mask;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire [31:0] tlSlaveXbar_out_0_a_bits_data;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_out_0_a_bits_corrupt;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_out_0_d_ready;	// src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_out_0_d_valid = tlSlaveXbar_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_out_0_d_bits_opcode = tlSlaveXbar_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_out_0_d_bits_size = tlSlaveXbar_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [4:0]  tlSlaveXbar__requestDOI_uncommonBits_T = tlSlaveXbar_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [31:0] tlSlaveXbar_out_0_d_bits_data = tlSlaveXbar_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_in_0_a_ready;	// src/main/scala/tilelink/Xbar.scala:155:18
  wire        slaveNodeOut_a_ready = tlSlaveXbar_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        slaveNodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlSlaveXbar_in_0_a_valid = tlSlaveXbar_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  slaveNodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  tlSlaveXbar_in_0_a_bits_opcode = tlSlaveXbar_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  slaveNodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  tlSlaveXbar_in_0_a_bits_param = tlSlaveXbar_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  slaveNodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  tlSlaveXbar_in_0_a_bits_size = tlSlaveXbar_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [4:0]  slaveNodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [4:0]  tlSlaveXbar_in_0_a_bits_source = tlSlaveXbar_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [31:0] slaveNodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] tlSlaveXbar__requestAIO_T = tlSlaveXbar_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [3:0]  slaveNodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  tlSlaveXbar_in_0_a_bits_mask = tlSlaveXbar_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [31:0] slaveNodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] tlSlaveXbar_in_0_a_bits_data = tlSlaveXbar_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire        slaveNodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlSlaveXbar_in_0_a_bits_corrupt = tlSlaveXbar_nodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire        slaveNodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlSlaveXbar_in_0_d_ready = tlSlaveXbar_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire        tlSlaveXbar_in_0_d_valid;	// src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  tlSlaveXbar_in_0_d_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:155:18
  wire        slaveNodeOut_d_valid = tlSlaveXbar_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  slaveNodeOut_d_bits_opcode = tlSlaveXbar_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlSlaveXbar_in_0_d_bits_size;	// src/main/scala/tilelink/Xbar.scala:155:18
  wire [4:0]  tlSlaveXbar_in_0_d_bits_source;	// src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  slaveNodeOut_d_bits_size = tlSlaveXbar_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [4:0]  slaveNodeOut_d_bits_source = tlSlaveXbar_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlSlaveXbar_in_0_d_bits_data;	// src/main/scala/tilelink/Xbar.scala:155:18
  wire [31:0] slaveNodeOut_d_bits_data = tlSlaveXbar_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlSlaveXbar_portsAOI_filtered_0_ready;	// src/main/scala/tilelink/Xbar.scala:348:24
  assign tlSlaveXbar_nodeIn_a_ready = tlSlaveXbar_in_0_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire        tlSlaveXbar_portsAOI_filtered_0_valid = tlSlaveXbar_in_0_a_valid;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [2:0]  tlSlaveXbar_portsAOI_filtered_0_bits_opcode =
    tlSlaveXbar_in_0_a_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [2:0]  tlSlaveXbar_portsAOI_filtered_0_bits_param = tlSlaveXbar_in_0_a_bits_param;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [2:0]  tlSlaveXbar_portsAOI_filtered_0_bits_size = tlSlaveXbar_in_0_a_bits_size;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [4:0]  tlSlaveXbar_portsAOI_filtered_0_bits_source =
    tlSlaveXbar_in_0_a_bits_source;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [31:0] tlSlaveXbar_portsAOI_filtered_0_bits_address = tlSlaveXbar__requestAIO_T;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [3:0]  tlSlaveXbar_portsAOI_filtered_0_bits_mask = tlSlaveXbar_in_0_a_bits_mask;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire [31:0] tlSlaveXbar_portsAOI_filtered_0_bits_data = tlSlaveXbar_in_0_a_bits_data;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire        tlSlaveXbar_portsAOI_filtered_0_bits_corrupt =
    tlSlaveXbar_in_0_a_bits_corrupt;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire        tlSlaveXbar_portsDIO_filtered_0_ready = tlSlaveXbar_in_0_d_ready;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire        tlSlaveXbar_portsDIO_filtered_0_valid;	// src/main/scala/tilelink/Xbar.scala:348:24
  assign tlSlaveXbar_nodeIn_d_valid = tlSlaveXbar_in_0_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  tlSlaveXbar_portsDIO_filtered_0_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:348:24
  assign tlSlaveXbar_nodeIn_d_bits_opcode = tlSlaveXbar_in_0_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [2:0]  tlSlaveXbar_portsDIO_filtered_0_bits_size;	// src/main/scala/tilelink/Xbar.scala:348:24
  assign tlSlaveXbar_nodeIn_d_bits_size = tlSlaveXbar_in_0_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [4:0]  tlSlaveXbar_portsDIO_filtered_0_bits_source;	// src/main/scala/tilelink/Xbar.scala:348:24
  assign tlSlaveXbar_nodeIn_d_bits_source = tlSlaveXbar_in_0_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  wire [31:0] tlSlaveXbar_portsDIO_filtered_0_bits_data;	// src/main/scala/tilelink/Xbar.scala:348:24
  assign tlSlaveXbar_nodeIn_d_bits_data = tlSlaveXbar_in_0_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17, src/main/scala/tilelink/Xbar.scala:155:18
  assign tlSlaveXbar_portsAOI_filtered_0_ready = tlSlaveXbar_out_0_a_ready;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  wire        tlSlaveXbar_nodeOut_a_valid = tlSlaveXbar_out_0_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_nodeOut_a_bits_opcode = tlSlaveXbar_out_0_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_nodeOut_a_bits_param = tlSlaveXbar_out_0_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [2:0]  tlSlaveXbar_nodeOut_a_bits_size = tlSlaveXbar_out_0_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [4:0]  tlSlaveXbar_nodeOut_a_bits_source = tlSlaveXbar_out_0_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [31:0] tlSlaveXbar_nodeOut_a_bits_address = tlSlaveXbar_out_0_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [3:0]  tlSlaveXbar_nodeOut_a_bits_mask = tlSlaveXbar_out_0_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire [31:0] tlSlaveXbar_nodeOut_a_bits_data = tlSlaveXbar_out_0_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_nodeOut_a_bits_corrupt = tlSlaveXbar_out_0_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  wire        tlSlaveXbar_nodeOut_d_ready = tlSlaveXbar_out_0_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Xbar.scala:212:19
  assign tlSlaveXbar_portsDIO_filtered_0_valid = tlSlaveXbar_out_0_d_valid;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_portsDIO_filtered_0_bits_opcode = tlSlaveXbar_out_0_d_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_portsDIO_filtered_0_bits_size = tlSlaveXbar_out_0_d_bits_size;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  wire [4:0]  tlSlaveXbar_requestDOI_uncommonBits =
    tlSlaveXbar__requestDOI_uncommonBits_T;	// src/main/scala/diplomacy/Parameters.scala:52:56, src/main/scala/tilelink/Xbar.scala:212:19
  assign tlSlaveXbar_portsDIO_filtered_0_bits_source =
    tlSlaveXbar__requestDOI_uncommonBits_T;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_portsDIO_filtered_0_bits_data = tlSlaveXbar_out_0_d_bits_data;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  wire [12:0] tlSlaveXbar__beatsAI_decode_T_1 = 13'h3F << tlSlaveXbar_in_0_a_bits_size;	// src/main/scala/tilelink/Xbar.scala:155:18, src/main/scala/util/package.scala:243:71
  wire [3:0]  tlSlaveXbar_beatsAI_decode = ~(tlSlaveXbar__beatsAI_decode_T_1[5:2]);	// src/main/scala/tilelink/Edges.scala:221:59, src/main/scala/util/package.scala:243:{46,71,76}
  wire        tlSlaveXbar_beatsAI_opdata = ~(tlSlaveXbar_in_0_a_bits_opcode[2]);	// src/main/scala/tilelink/Edges.scala:93:{28,37}, src/main/scala/tilelink/Xbar.scala:155:18
  wire [3:0]  tlSlaveXbar_beatsAI_0 =
    tlSlaveXbar_beatsAI_opdata ? tlSlaveXbar_beatsAI_decode : 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Edges.scala:93:28, :221:59, :222:14
  wire [12:0] tlSlaveXbar__beatsDO_decode_T_1 = 13'h3F << tlSlaveXbar_out_0_d_bits_size;	// src/main/scala/tilelink/Xbar.scala:212:19, src/main/scala/util/package.scala:243:71
  wire [3:0]  tlSlaveXbar_beatsDO_decode = ~(tlSlaveXbar__beatsDO_decode_T_1[5:2]);	// src/main/scala/tilelink/Edges.scala:221:59, src/main/scala/util/package.scala:243:{46,71,76}
  wire        tlSlaveXbar_beatsDO_opdata = tlSlaveXbar_out_0_d_bits_opcode[0];	// src/main/scala/tilelink/Edges.scala:107:36, src/main/scala/tilelink/Xbar.scala:212:19
  wire [3:0]  tlSlaveXbar_beatsDO_0 =
    tlSlaveXbar_beatsDO_opdata ? tlSlaveXbar_beatsDO_decode : 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, src/main/scala/tilelink/Edges.scala:107:36, :221:59, :222:14
  assign tlSlaveXbar_in_0_a_ready = tlSlaveXbar_portsAOI_filtered_0_ready;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  assign tlSlaveXbar_out_0_a_valid = tlSlaveXbar_portsAOI_filtered_0_valid;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_opcode = tlSlaveXbar_portsAOI_filtered_0_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_param = tlSlaveXbar_portsAOI_filtered_0_bits_param;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_size = tlSlaveXbar_portsAOI_filtered_0_bits_size;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_source = tlSlaveXbar_portsAOI_filtered_0_bits_source;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_address = tlSlaveXbar_portsAOI_filtered_0_bits_address;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_mask = tlSlaveXbar_portsAOI_filtered_0_bits_mask;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_data = tlSlaveXbar_portsAOI_filtered_0_bits_data;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_a_bits_corrupt = tlSlaveXbar_portsAOI_filtered_0_bits_corrupt;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_out_0_d_ready = tlSlaveXbar_portsDIO_filtered_0_ready;	// src/main/scala/tilelink/Xbar.scala:212:19, :348:24
  assign tlSlaveXbar_in_0_d_valid = tlSlaveXbar_portsDIO_filtered_0_valid;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  assign tlSlaveXbar_in_0_d_bits_opcode = tlSlaveXbar_portsDIO_filtered_0_bits_opcode;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  assign tlSlaveXbar_in_0_d_bits_size = tlSlaveXbar_portsDIO_filtered_0_bits_size;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  assign tlSlaveXbar_in_0_d_bits_source = tlSlaveXbar_portsDIO_filtered_0_bits_source;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  assign tlSlaveXbar_in_0_d_bits_data = tlSlaveXbar_portsDIO_filtered_0_bits_data;	// src/main/scala/tilelink/Xbar.scala:155:18, :348:24
  wire        hartidOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_nodeIn;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_nodeOut = broadcast_nodeIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        broadcast_x1_nodeOut = broadcast_nodeIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        hartIdSinkNodeIn = broadcast_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        traceSourceNodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeOut_insns_0_valid = broadcast_3_nodeIn_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] traceSourceNodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_nodeOut_insns_0_iaddr = broadcast_3_nodeIn_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] traceSourceNodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_nodeOut_insns_0_insn = broadcast_3_nodeIn_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  traceSourceNodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  broadcast_3_nodeOut_insns_0_priv = broadcast_3_nodeIn_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        traceSourceNodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeOut_insns_0_exception =
    broadcast_3_nodeIn_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        traceSourceNodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeOut_insns_0_interrupt =
    broadcast_3_nodeIn_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] traceSourceNodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_nodeOut_insns_0_cause = broadcast_3_nodeIn_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] traceSourceNodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_nodeOut_insns_0_tval = broadcast_3_nodeIn_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [63:0] traceSourceNodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_nodeOut_time = broadcast_3_nodeIn_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        bpwatchSourceNodeOut_0_valid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  bpwatchSourceNodeOut_0_action;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeIn_a_ready = widget_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_valid = widget_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  widget_nodeIn_d_bits_opcode = widget_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [1:0]  widget_nodeIn_d_bits_param = widget_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  widget_nodeIn_d_bits_size = widget_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeIn_d_bits_sink = widget_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeIn_d_bits_denied = widget_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] widget_nodeIn_d_bits_data = widget_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeIn_d_bits_corrupt = widget_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_a_valid = widget_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  widget_nodeOut_a_bits_opcode = widget_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  widget_nodeOut_a_bits_param = widget_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  widget_nodeOut_a_bits_size = widget_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] widget_nodeOut_a_bits_address = widget_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_a_bits_user_amba_prot_bufferable =
    widget_nodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_a_bits_user_amba_prot_modifiable =
    widget_nodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_a_bits_user_amba_prot_readalloc =
    widget_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_a_bits_user_amba_prot_writealloc =
    widget_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_a_bits_user_amba_prot_privileged =
    widget_nodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  widget_nodeOut_a_bits_mask = widget_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] widget_nodeOut_a_bits_data = widget_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_nodeOut_d_ready = widget_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeIn_a_ready = widget_1_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_1_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_d_valid = widget_1_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  widget_1_nodeIn_d_bits_opcode = widget_1_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [1:0]  widget_1_nodeIn_d_bits_param = widget_1_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  widget_1_nodeIn_d_bits_size = widget_1_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeIn_d_bits_sink = widget_1_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeIn_d_bits_denied = widget_1_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] widget_1_nodeIn_d_bits_data = widget_1_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeIn_d_bits_corrupt = widget_1_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeOut_a_valid = widget_1_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] widget_1_nodeOut_a_bits_address = widget_1_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_readalloc =
    widget_1_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_writealloc =
    widget_1_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_nodeIn_a_ready = buffer_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  buffer_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] buffer_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  buffer_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] buffer_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_nodeIn_d_valid = buffer_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  buffer_nodeIn_d_bits_opcode = buffer_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [1:0]  buffer_nodeIn_d_bits_param = buffer_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  buffer_nodeIn_d_bits_size = buffer_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_nodeIn_d_bits_source = buffer_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_nodeIn_d_bits_sink = buffer_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_nodeIn_d_bits_denied = buffer_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] buffer_nodeIn_d_bits_data = buffer_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_nodeIn_d_bits_corrupt = buffer_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_a_ready = buffer_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_valid = buffer_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlOtherMastersNodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_a_bits_opcode = buffer_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlOtherMastersNodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_a_bits_param = buffer_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  tlOtherMastersNodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_a_bits_size = buffer_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_source = buffer_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlOtherMastersNodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeOut_a_bits_address = buffer_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  tlOtherMastersNodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_a_bits_mask = buffer_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlOtherMastersNodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeOut_a_bits_data = buffer_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_ready = buffer_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_d_valid = buffer_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlOtherMastersNodeOut_d_bits_opcode = buffer_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [1:0]  tlOtherMastersNodeOut_d_bits_param = buffer_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  tlOtherMastersNodeOut_d_bits_size = buffer_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_d_bits_source = buffer_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_d_bits_sink = buffer_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_d_bits_denied = buffer_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlOtherMastersNodeOut_d_bits_data = buffer_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeOut_d_bits_corrupt = buffer_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        slaveNodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_1_nodeIn_a_ready = buffer_1_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        slaveNodeIn_a_valid = buffer_1_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  slaveNodeIn_a_bits_opcode = buffer_1_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  slaveNodeIn_a_bits_param = buffer_1_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  slaveNodeIn_a_bits_size = buffer_1_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [4:0]  slaveNodeIn_a_bits_source = buffer_1_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] slaveNodeIn_a_bits_address = buffer_1_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  slaveNodeIn_a_bits_mask = buffer_1_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] slaveNodeIn_a_bits_data = buffer_1_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        slaveNodeIn_a_bits_corrupt = buffer_1_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        slaveNodeIn_d_ready = buffer_1_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        slaveNodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_1_nodeIn_d_valid = buffer_1_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  slaveNodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_1_nodeIn_d_bits_opcode = buffer_1_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  slaveNodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_1_nodeIn_d_bits_size = buffer_1_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [4:0]  slaveNodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [4:0]  buffer_1_nodeIn_d_bits_source = buffer_1_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] slaveNodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] buffer_1_nodeIn_d_bits_data = buffer_1_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_valid = buffer_1_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_opcode = buffer_1_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_param = buffer_1_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_size = buffer_1_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_source = buffer_1_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_address = buffer_1_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_mask = buffer_1_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_data = buffer_1_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_bits_corrupt = buffer_1_nodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_d_ready = buffer_1_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_a_ready = tlOtherMastersNodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_valid = tlOtherMastersNodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlOtherMastersNodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_opcode = tlOtherMastersNodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlOtherMastersNodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_param = tlOtherMastersNodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  tlOtherMastersNodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_size = tlOtherMastersNodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_source = tlOtherMastersNodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlOtherMastersNodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_address = tlOtherMastersNodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  tlOtherMastersNodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_mask = tlOtherMastersNodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlOtherMastersNodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_a_bits_data = tlOtherMastersNodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeIn_d_ready = tlOtherMastersNodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_d_valid = tlOtherMastersNodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  tlOtherMastersNodeIn_d_bits_opcode = tlOtherMastersNodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [1:0]  tlOtherMastersNodeIn_d_bits_param = tlOtherMastersNodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [3:0]  tlOtherMastersNodeIn_d_bits_size = tlOtherMastersNodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_d_bits_source = tlOtherMastersNodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_d_bits_sink = tlOtherMastersNodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_d_bits_denied = tlOtherMastersNodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [31:0] tlOtherMastersNodeIn_d_bits_data = tlOtherMastersNodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        tlOtherMastersNodeIn_d_bits_corrupt = tlOtherMastersNodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_valid = tlOtherMastersNodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_opcode = tlOtherMastersNodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_param = tlOtherMastersNodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_size = tlOtherMastersNodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_source = tlOtherMastersNodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_address = tlOtherMastersNodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_mask = tlOtherMastersNodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_data = tlOtherMastersNodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_d_ready = tlOtherMastersNodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_nodeIn = hartidOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign hartidOut = hartidIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_valid = traceSourceNodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_iaddr = traceSourceNodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_insn = traceSourceNodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_priv = traceSourceNodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_exception = traceSourceNodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_interrupt = traceSourceNodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_cause = traceSourceNodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_insns_0_tval = traceSourceNodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeIn_time = traceSourceNodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        broadcast_4_nodeIn_0_valid_0 = bpwatchSourceNodeOut_0_valid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire [2:0]  broadcast_4_nodeIn_0_action = bpwatchSourceNodeOut_0_action;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        int_localOut_0 = int_localIn_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        x1_int_localOut_0 = x1_int_localIn_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        x1_int_localOut_1 = x1_int_localIn_1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        x1_int_localOut_1_0 = x1_int_localIn_1_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeIn_a_ready = slaveNodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_valid = slaveNodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_opcode = slaveNodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_param = slaveNodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_size = slaveNodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_source = slaveNodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_address = slaveNodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_mask = slaveNodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_data = slaveNodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_a_bits_corrupt = slaveNodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlSlaveXbar_nodeIn_d_ready = slaveNodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeIn_d_valid = slaveNodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeIn_d_bits_opcode = slaveNodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeIn_d_bits_size = slaveNodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeIn_d_bits_source = slaveNodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeIn_d_bits_data = slaveNodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_a_ready = slaveNodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_valid = slaveNodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_opcode = slaveNodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_param = slaveNodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_size = slaveNodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_source = slaveNodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_address = slaveNodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_mask = slaveNodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_data = slaveNodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_a_bits_corrupt = slaveNodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign slaveNodeOut_d_ready = slaveNodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_d_valid = slaveNodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_d_bits_opcode = slaveNodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_d_bits_size = slaveNodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_d_bits_source = slaveNodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_1_nodeOut_d_bits_data = slaveNodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  reg         wfiNodeOut_0_REG;	// src/main/scala/tile/Interrupts.scala:126:36
  wire        wfiNodeOut_0 = wfiNodeOut_0_REG;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/Interrupts.scala:126:36
  always @(posedge clock) begin
    if (reset)
      wfiNodeOut_0_REG <= 1'h0;	// src/main/scala/diplomacy/LazyModule.scala:374:18, src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17, src/main/scala/rocket/Frontend.scala:386:28, src/main/scala/rocket/HellaCache.scala:269:43, :286:25, src/main/scala/rocket/PTW.scala:801:19, src/main/scala/tile/BaseTile.scala:218:42, :294:19, src/main/scala/tile/Interrupts.scala:126:36, src/main/scala/tile/RocketTile.scala:60:15, :127:20, src/main/scala/tilelink/Edges.scala:103:36, src/main/scala/tilelink/Fragmenter.scala:335:34, src/main/scala/tilelink/Xbar.scala:155:18, :212:19, :348:24
    else
      wfiNodeOut_0_REG <= _core_io_wfi;	// src/main/scala/tile/Interrupts.scala:126:36, src/main/scala/tile/RocketTile.scala:127:20
  end // always @(posedge)
  wire tlMasterXbar_clock;
    wire tlMasterXbar_reset;
    wire tlMasterXbar_auto_in_1_a_ready;
    wire tlMasterXbar_auto_in_1_a_valid;
    wire[31:0] tlMasterXbar_auto_in_1_a_bits_address;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_in_1_d_valid;
    wire[2:0] tlMasterXbar_auto_in_1_d_bits_opcode;
    wire[1:0] tlMasterXbar_auto_in_1_d_bits_param;
    wire[3:0] tlMasterXbar_auto_in_1_d_bits_size;
    wire tlMasterXbar_auto_in_1_d_bits_sink;
    wire tlMasterXbar_auto_in_1_d_bits_denied;
    wire[31:0] tlMasterXbar_auto_in_1_d_bits_data;
    wire tlMasterXbar_auto_in_1_d_bits_corrupt;
    wire tlMasterXbar_auto_in_0_a_ready;
    wire tlMasterXbar_auto_in_0_a_valid;
    wire[2:0] tlMasterXbar_auto_in_0_a_bits_opcode;
    wire[2:0] tlMasterXbar_auto_in_0_a_bits_param;
    wire[3:0] tlMasterXbar_auto_in_0_a_bits_size;
    wire[31:0] tlMasterXbar_auto_in_0_a_bits_address;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_privileged;
    wire[3:0] tlMasterXbar_auto_in_0_a_bits_mask;
    wire[31:0] tlMasterXbar_auto_in_0_a_bits_data;
    wire tlMasterXbar_auto_in_0_d_ready;
    wire tlMasterXbar_auto_in_0_d_valid;
    wire[2:0] tlMasterXbar_auto_in_0_d_bits_opcode;
    wire[1:0] tlMasterXbar_auto_in_0_d_bits_param;
    wire[3:0] tlMasterXbar_auto_in_0_d_bits_size;
    wire tlMasterXbar_auto_in_0_d_bits_sink;
    wire tlMasterXbar_auto_in_0_d_bits_denied;
    wire[31:0] tlMasterXbar_auto_in_0_d_bits_data;
    wire tlMasterXbar_auto_in_0_d_bits_corrupt;
    wire tlMasterXbar_auto_out_a_ready;
    wire tlMasterXbar_auto_out_a_valid;
    wire[2:0] tlMasterXbar_auto_out_a_bits_opcode;
    wire[2:0] tlMasterXbar_auto_out_a_bits_param;
    wire[3:0] tlMasterXbar_auto_out_a_bits_size;
    wire tlMasterXbar_auto_out_a_bits_source;
    wire[31:0] tlMasterXbar_auto_out_a_bits_address;
    wire[3:0] tlMasterXbar_auto_out_a_bits_mask;
    wire[31:0] tlMasterXbar_auto_out_a_bits_data;
    wire tlMasterXbar_auto_out_d_ready;
    wire tlMasterXbar_auto_out_d_valid;
    wire[2:0] tlMasterXbar_auto_out_d_bits_opcode;
    wire[1:0] tlMasterXbar_auto_out_d_bits_param;
    wire[3:0] tlMasterXbar_auto_out_d_bits_size;
    wire tlMasterXbar_auto_out_d_bits_source;
    wire tlMasterXbar_auto_out_d_bits_sink;
    wire tlMasterXbar_auto_out_d_bits_denied;
    wire[31:0] tlMasterXbar_auto_out_d_bits_data;
    wire tlMasterXbar_auto_out_d_bits_corrupt;

    wire tlMasterXbar_nodeIn_a_valid = tlMasterXbar_auto_in_0_a_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_a_bits_opcode = tlMasterXbar_auto_in_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeIn_a_bits_param = tlMasterXbar_auto_in_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_a_bits_size = tlMasterXbar_auto_in_0_a_bits_size ; 
    wire[31:0] tlMasterXbar_nodeIn_a_bits_address = tlMasterXbar_auto_in_0_a_bits_address ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_bufferable = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_modifiable = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_readalloc = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_writealloc = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_privileged = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_privileged ; 
    wire[3:0] tlMasterXbar_nodeIn_a_bits_mask = tlMasterXbar_auto_in_0_a_bits_mask ; 
    wire[31:0] tlMasterXbar_nodeIn_a_bits_data = tlMasterXbar_auto_in_0_a_bits_data ; 
    wire tlMasterXbar_nodeIn_d_ready = tlMasterXbar_auto_in_0_d_ready ; 
    wire tlMasterXbar_nodeIn_1_a_valid = tlMasterXbar_auto_in_1_a_valid ; 
    wire[31:0] tlMasterXbar_nodeIn_1_a_bits_address = tlMasterXbar_auto_in_1_a_bits_address ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_readalloc = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_writealloc = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeOut_a_ready = tlMasterXbar_auto_out_a_ready ; 
    wire tlMasterXbar_nodeOut_d_valid = tlMasterXbar_auto_out_d_valid ; 
    wire[2:0] tlMasterXbar_nodeOut_d_bits_opcode = tlMasterXbar_auto_out_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_nodeOut_d_bits_param = tlMasterXbar_auto_out_d_bits_param ; 
    wire[3:0] tlMasterXbar_nodeOut_d_bits_size = tlMasterXbar_auto_out_d_bits_size ; 
    wire tlMasterXbar_nodeOut_d_bits_source = tlMasterXbar_auto_out_d_bits_source ; 
    wire tlMasterXbar_nodeOut_d_bits_sink = tlMasterXbar_auto_out_d_bits_sink ; 
    wire tlMasterXbar_nodeOut_d_bits_denied = tlMasterXbar_auto_out_d_bits_denied ; 
    wire[31:0] tlMasterXbar_nodeOut_d_bits_data = tlMasterXbar_auto_out_d_bits_data ; 
    wire tlMasterXbar_nodeOut_d_bits_corrupt = tlMasterXbar_auto_out_d_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_a_bits_source =1'h0; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_nodeIn_a_bits_corrupt =1'h0; 
    wire tlMasterXbar_nodeIn_d_bits_source =1'h0; 
    wire tlMasterXbar_nodeIn_1_a_bits_source =1'h0; 
    wire tlMasterXbar_nodeIn_1_a_bits_corrupt =1'h0; 
    wire tlMasterXbar_nodeIn_1_d_bits_source =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_nodeOut_a_bits_corrupt =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_in_0_a_bits_corrupt =1'h0; 
    wire tlMasterXbar_in_1_a_bits_source =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_in_1_a_bits_corrupt =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_out_0_a_bits_corrupt =1'h0; 
    wire tlMasterXbar_requestBOI_0_0 =1'h0; 
    wire tlMasterXbar_beatsAI_opdata_1 =1'h0; 
    wire tlMasterXbar_beatsCI_opdata =1'h0; 
    wire tlMasterXbar_beatsCI_opdata_1 =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_corrupt =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_source =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_corrupt =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_0_ready =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_0_valid =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_0_bits_source =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_0_bits_corrupt =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_1_ready =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_1_valid =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_1_bits_source =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_1_bits_corrupt =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_ready =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_valid =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_source =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_corrupt =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_ready =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_valid =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_source =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_corrupt =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_0_ready =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_0_valid =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_0_bits_sink =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_1_0_ready =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_1_0_valid =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_1_0_bits_sink =1'h0; 
    wire[1:0] tlMasterXbar_portsBIO_filtered_0_bits_param =2'h0; 
    wire[1:0] tlMasterXbar_portsBIO_filtered_1_bits_param =2'h0; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_secure =1'h1; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_bufferable =1'h1; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_modifiable =1'h1; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_privileged =1'h1; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_secure =1'h1; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_fetch =1'h1; 
    wire tlMasterXbar_nodeIn_1_d_ready =1'h1; 
    wire tlMasterXbar_in_0_a_bits_source =1'h1; 
    wire tlMasterXbar_in_1_d_ready =1'h1; 
    wire tlMasterXbar_requestAIO_0_0 =1'h1; 
    wire tlMasterXbar_requestAIO_1_0 =1'h1; 
    wire tlMasterXbar_requestCIO_0_0 =1'h1; 
    wire tlMasterXbar_requestCIO_1_0 =1'h1; 
    wire tlMasterXbar_requestBOI_0_1 =1'h1; 
    wire tlMasterXbar_beatsBO_opdata =1'h1; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_source =1'h1; 
    wire tlMasterXbar_portsDIO_filtered_1_ready =1'h1; 
    wire[2:0] tlMasterXbar_nodeIn_1_a_bits_opcode =3'h4; 
    wire[2:0] tlMasterXbar_in_1_a_bits_opcode =3'h4; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_1_0_bits_opcode =3'h4; 
    wire[2:0] tlMasterXbar_nodeIn_1_a_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_in_1_a_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_1_0_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_portsBIO_filtered_0_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_portsBIO_filtered_1_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_0_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_0_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_1_0_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_1_0_bits_param =3'h0; 
    wire[3:0] tlMasterXbar_nodeIn_1_a_bits_size =4'h6; 
    wire[3:0] tlMasterXbar_in_1_a_bits_size =4'h6; 
    wire[3:0] tlMasterXbar_portsAOI_filtered_1_0_bits_size =4'h6; 
    wire[3:0] tlMasterXbar_nodeIn_1_a_bits_mask =4'hF; 
    wire[3:0] tlMasterXbar_in_1_a_bits_mask =4'hF; 
    wire[3:0] tlMasterXbar_portsAOI_filtered_1_0_bits_mask =4'hF; 
    wire[31:0] tlMasterXbar_nodeIn_1_a_bits_data =32'h0; 
    wire[31:0] tlMasterXbar_in_1_a_bits_data =32'h0; 
    wire[31:0] tlMasterXbar_portsAOI_filtered_1_0_bits_data =32'h0; 
    wire[31:0] tlMasterXbar_portsBIO_filtered_0_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_portsBIO_filtered_0_bits_data =32'h0; 
    wire[31:0] tlMasterXbar_portsBIO_filtered_1_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_portsBIO_filtered_1_bits_data =32'h0; 
    wire[31:0] tlMasterXbar_portsCOI_filtered_0_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_portsCOI_filtered_0_bits_data =32'h0; 
    wire[31:0] tlMasterXbar_portsCOI_filtered_1_0_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_portsCOI_filtered_1_0_bits_data =32'h0; 
    wire[9:0] tlMasterXbar_beatsAI_1 =10'h0; 
    wire[9:0] tlMasterXbar_beatsBO_decode =10'h0; 
    wire[9:0] tlMasterXbar_beatsBO_0 =10'h0; 
    wire[9:0] tlMasterXbar_beatsCI_decode =10'h0; 
    wire[9:0] tlMasterXbar_beatsCI_0 =10'h0; 
    wire[9:0] tlMasterXbar_beatsCI_decode_1 =10'h0; 
    wire[9:0] tlMasterXbar_beatsCI_1 =10'h0; 
    wire[9:0] tlMasterXbar_maskedBeats_1 =10'h0; 
    wire[9:0] tlMasterXbar_beatsAI_decode_1 =10'hF; 
    wire[3:0] tlMasterXbar_portsBIO_filtered_0_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_portsBIO_filtered_0_bits_mask =4'h0; 
    wire[3:0] tlMasterXbar_portsBIO_filtered_1_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_portsBIO_filtered_1_bits_mask =4'h0; 
    wire[3:0] tlMasterXbar_portsCOI_filtered_0_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_portsCOI_filtered_1_0_bits_size =4'h0; 
    wire tlMasterXbar_in_0_a_ready ; 
    wire tlMasterXbar_in_0_a_valid = tlMasterXbar_nodeIn_a_valid ; 
    wire[2:0] tlMasterXbar_in_0_a_bits_opcode = tlMasterXbar_nodeIn_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_in_0_a_bits_param = tlMasterXbar_nodeIn_a_bits_param ; 
    wire[3:0] tlMasterXbar_in_0_a_bits_size = tlMasterXbar_nodeIn_a_bits_size ; 
    wire[31:0] tlMasterXbar_in_0_a_bits_address = tlMasterXbar_nodeIn_a_bits_address ; 
    wire[3:0] tlMasterXbar_in_0_a_bits_mask = tlMasterXbar_nodeIn_a_bits_mask ; 
    wire[31:0] tlMasterXbar_in_0_a_bits_data = tlMasterXbar_nodeIn_a_bits_data ; 
    wire tlMasterXbar_in_0_d_ready = tlMasterXbar_nodeIn_d_ready ; 
    wire tlMasterXbar_in_0_d_valid ; 
    wire[2:0] tlMasterXbar_in_0_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_in_0_d_bits_param ; 
    wire[3:0] tlMasterXbar_in_0_d_bits_size ; 
    wire tlMasterXbar_in_0_d_bits_sink ; 
    wire tlMasterXbar_in_0_d_bits_denied ; 
    wire[31:0] tlMasterXbar_in_0_d_bits_data ; 
    wire tlMasterXbar_in_0_d_bits_corrupt ; 
    wire tlMasterXbar_in_1_a_ready ; 
    wire tlMasterXbar_in_1_a_valid = tlMasterXbar_nodeIn_1_a_valid ; 
    wire[31:0] tlMasterXbar_in_1_a_bits_address = tlMasterXbar_nodeIn_1_a_bits_address ; 
    wire tlMasterXbar_in_1_d_valid ; 
    wire[2:0] tlMasterXbar_in_1_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_in_1_d_bits_param ; 
    wire[3:0] tlMasterXbar_in_1_d_bits_size ; 
    wire tlMasterXbar_in_1_d_bits_sink ; 
    wire tlMasterXbar_in_1_d_bits_denied ; 
    wire[31:0] tlMasterXbar_in_1_d_bits_data ; 
    wire tlMasterXbar_in_1_d_bits_corrupt ; 
    wire tlMasterXbar_out_0_a_ready = tlMasterXbar_nodeOut_a_ready ; 
    wire tlMasterXbar_out_0_a_valid ; 
    wire[2:0] tlMasterXbar_out_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_out_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_out_0_a_bits_size ; 
    wire tlMasterXbar_out_0_a_bits_source ; 
    wire[31:0] tlMasterXbar_out_0_a_bits_address ; 
    wire[3:0] tlMasterXbar_out_0_a_bits_mask ; 
    wire[31:0] tlMasterXbar_out_0_a_bits_data ; 
    wire tlMasterXbar_out_0_d_ready ; 
    wire tlMasterXbar_out_0_d_valid = tlMasterXbar_nodeOut_d_valid ; 
    wire[2:0] tlMasterXbar_out_0_d_bits_opcode = tlMasterXbar_nodeOut_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_out_0_d_bits_param = tlMasterXbar_nodeOut_d_bits_param ; 
    wire[3:0] tlMasterXbar_out_0_d_bits_size = tlMasterXbar_nodeOut_d_bits_size ; 
    wire tlMasterXbar_out_0_d_bits_source = tlMasterXbar_nodeOut_d_bits_source ; 
    wire tlMasterXbar_out_0_d_bits_sink = tlMasterXbar_nodeOut_d_bits_sink ; 
    wire tlMasterXbar_out_0_d_bits_denied = tlMasterXbar_nodeOut_d_bits_denied ; 
    wire[31:0] tlMasterXbar_out_0_d_bits_data = tlMasterXbar_nodeOut_d_bits_data ; 
    wire tlMasterXbar_out_0_d_bits_corrupt = tlMasterXbar_nodeOut_d_bits_corrupt ; 
    wire tlMasterXbar_portsAOI_filtered_0_ready ; 
    wire tlMasterXbar_nodeIn_a_ready = tlMasterXbar_in_0_a_ready ; 
    wire tlMasterXbar_portsAOI_filtered_0_valid = tlMasterXbar_in_0_a_valid ; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_0_bits_opcode = tlMasterXbar_in_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_0_bits_param = tlMasterXbar_in_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_portsAOI_filtered_0_bits_size = tlMasterXbar_in_0_a_bits_size ; 
    wire[31:0] tlMasterXbar_portsAOI_filtered_0_bits_address = tlMasterXbar_in_0_a_bits_address ; 
    wire[3:0] tlMasterXbar_portsAOI_filtered_0_bits_mask = tlMasterXbar_in_0_a_bits_mask ; 
    wire[31:0] tlMasterXbar_portsAOI_filtered_0_bits_data = tlMasterXbar_in_0_a_bits_data ; 
    wire tlMasterXbar_portsDIO_filtered_0_ready = tlMasterXbar_in_0_d_ready ; 
    wire tlMasterXbar_portsDIO_filtered_0_valid ; 
    wire tlMasterXbar_nodeIn_d_valid = tlMasterXbar_in_0_d_valid ; 
    wire[2:0] tlMasterXbar_portsDIO_filtered_0_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeIn_d_bits_opcode = tlMasterXbar_in_0_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_0_bits_param ; 
    wire[1:0] tlMasterXbar_nodeIn_d_bits_param = tlMasterXbar_in_0_d_bits_param ; 
    wire[3:0] tlMasterXbar_portsDIO_filtered_0_bits_size ; 
    wire[3:0] tlMasterXbar_nodeIn_d_bits_size = tlMasterXbar_in_0_d_bits_size ; 
    wire tlMasterXbar_portsDIO_filtered_0_bits_source ; 
    wire tlMasterXbar_portsDIO_filtered_0_bits_sink ; 
    wire tlMasterXbar_nodeIn_d_bits_sink = tlMasterXbar_in_0_d_bits_sink ; 
    wire tlMasterXbar_portsDIO_filtered_0_bits_denied ; 
    wire tlMasterXbar_nodeIn_d_bits_denied = tlMasterXbar_in_0_d_bits_denied ; 
    wire[31:0] tlMasterXbar_portsDIO_filtered_0_bits_data ; 
    wire[31:0] tlMasterXbar_nodeIn_d_bits_data = tlMasterXbar_in_0_d_bits_data ; 
    wire tlMasterXbar_portsDIO_filtered_0_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_d_bits_corrupt = tlMasterXbar_in_0_d_bits_corrupt ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_ready ; 
    wire tlMasterXbar_nodeIn_1_a_ready = tlMasterXbar_in_1_a_ready ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_valid = tlMasterXbar_in_1_a_valid ; 
    wire[31:0] tlMasterXbar_portsAOI_filtered_1_0_bits_address = tlMasterXbar_in_1_a_bits_address ; 
    wire tlMasterXbar_portsDIO_filtered_1_valid ; 
    wire tlMasterXbar_nodeIn_1_d_valid = tlMasterXbar_in_1_d_valid ; 
    wire[2:0] tlMasterXbar_portsDIO_filtered_1_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeIn_1_d_bits_opcode = tlMasterXbar_in_1_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_1_bits_param ; 
    wire[1:0] tlMasterXbar_nodeIn_1_d_bits_param = tlMasterXbar_in_1_d_bits_param ; 
    wire[3:0] tlMasterXbar_portsDIO_filtered_1_bits_size ; 
    wire[3:0] tlMasterXbar_nodeIn_1_d_bits_size = tlMasterXbar_in_1_d_bits_size ; 
    wire tlMasterXbar_portsDIO_filtered_1_bits_source ; 
    wire tlMasterXbar_portsDIO_filtered_1_bits_sink ; 
    wire tlMasterXbar_nodeIn_1_d_bits_sink = tlMasterXbar_in_1_d_bits_sink ; 
    wire tlMasterXbar_portsDIO_filtered_1_bits_denied ; 
    wire tlMasterXbar_nodeIn_1_d_bits_denied = tlMasterXbar_in_1_d_bits_denied ; 
    wire[31:0] tlMasterXbar_portsDIO_filtered_1_bits_data ; 
    wire[31:0] tlMasterXbar_nodeIn_1_d_bits_data = tlMasterXbar_in_1_d_bits_data ; 
    wire tlMasterXbar_portsDIO_filtered_1_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_1_d_bits_corrupt = tlMasterXbar_in_1_d_bits_corrupt ; 
    wire tlMasterXbar_nodeOut_a_valid = tlMasterXbar_out_0_a_valid ; 
    wire[2:0] tlMasterXbar_nodeOut_a_bits_opcode = tlMasterXbar_out_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeOut_a_bits_param = tlMasterXbar_out_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_nodeOut_a_bits_size = tlMasterXbar_out_0_a_bits_size ; 
    wire tlMasterXbar_muxState_0 ; 
    wire tlMasterXbar_nodeOut_a_bits_source = tlMasterXbar_out_0_a_bits_source ; 
    wire[31:0] tlMasterXbar_nodeOut_a_bits_address = tlMasterXbar_out_0_a_bits_address ; 
    wire[3:0] tlMasterXbar_nodeOut_a_bits_mask = tlMasterXbar_out_0_a_bits_mask ; 
    wire[31:0] tlMasterXbar_nodeOut_a_bits_data = tlMasterXbar_out_0_a_bits_data ; 
    wire tlMasterXbar_nodeOut_d_ready = tlMasterXbar_out_0_d_ready ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_opcode = tlMasterXbar_out_0_d_bits_opcode ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_opcode = tlMasterXbar_out_0_d_bits_opcode ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_param = tlMasterXbar_out_0_d_bits_param ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_param = tlMasterXbar_out_0_d_bits_param ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_size = tlMasterXbar_out_0_d_bits_size ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_size = tlMasterXbar_out_0_d_bits_size ; 
    wire tlMasterXbar_requestDOI_0_0 = tlMasterXbar_out_0_d_bits_source ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_source = tlMasterXbar_out_0_d_bits_source ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_source = tlMasterXbar_out_0_d_bits_source ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_sink = tlMasterXbar_out_0_d_bits_sink ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_sink = tlMasterXbar_out_0_d_bits_sink ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_denied = tlMasterXbar_out_0_d_bits_denied ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_denied = tlMasterXbar_out_0_d_bits_denied ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_data = tlMasterXbar_out_0_d_bits_data ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_data = tlMasterXbar_out_0_d_bits_data ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_corrupt = tlMasterXbar_out_0_d_bits_corrupt ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_corrupt = tlMasterXbar_out_0_d_bits_corrupt ; 
    wire tlMasterXbar_requestDOI_0_1 =~ tlMasterXbar_out_0_d_bits_source ; 
    wire[26:0] tlMasterXbar__beatsAI_decode_T_1 =27'hFFF<< tlMasterXbar_in_0_a_bits_size ; 
    wire[9:0] tlMasterXbar_beatsAI_decode =~( tlMasterXbar__beatsAI_decode_T_1 [11:2]); 
    wire tlMasterXbar_beatsAI_opdata =~( tlMasterXbar_in_0_a_bits_opcode [2]); 
    wire[9:0] tlMasterXbar_beatsAI_0 = tlMasterXbar_beatsAI_opdata  ?  tlMasterXbar_beatsAI_decode :10'h0; 
    wire[26:0] tlMasterXbar__beatsDO_decode_T_1 =27'hFFF<< tlMasterXbar_out_0_d_bits_size ; 
    wire[9:0] tlMasterXbar_beatsDO_decode =~( tlMasterXbar__beatsDO_decode_T_1 [11:2]); 
    wire tlMasterXbar_beatsDO_opdata = tlMasterXbar_out_0_d_bits_opcode [0]; 
    wire[9:0] tlMasterXbar_beatsDO_0 = tlMasterXbar_beatsDO_opdata  ?  tlMasterXbar_beatsDO_decode :10'h0; 
  assign  tlMasterXbar_in_0_a_ready = tlMasterXbar_portsAOI_filtered_0_ready ; 
  assign  tlMasterXbar_in_1_a_ready = tlMasterXbar_portsAOI_filtered_1_0_ready ; 
  assign  tlMasterXbar_in_0_d_valid = tlMasterXbar_portsDIO_filtered_0_valid ; 
  assign  tlMasterXbar_in_0_d_bits_opcode = tlMasterXbar_portsDIO_filtered_0_bits_opcode ; 
  assign  tlMasterXbar_in_0_d_bits_param = tlMasterXbar_portsDIO_filtered_0_bits_param ; 
  assign  tlMasterXbar_in_0_d_bits_size = tlMasterXbar_portsDIO_filtered_0_bits_size ; 
    wire tlMasterXbar_in_0_d_bits_source = tlMasterXbar_portsDIO_filtered_0_bits_source ; 
  assign  tlMasterXbar_in_0_d_bits_sink = tlMasterXbar_portsDIO_filtered_0_bits_sink ; 
  assign  tlMasterXbar_in_0_d_bits_denied = tlMasterXbar_portsDIO_filtered_0_bits_denied ; 
  assign  tlMasterXbar_in_0_d_bits_data = tlMasterXbar_portsDIO_filtered_0_bits_data ; 
  assign  tlMasterXbar_in_0_d_bits_corrupt = tlMasterXbar_portsDIO_filtered_0_bits_corrupt ; 
  assign  tlMasterXbar_in_1_d_valid = tlMasterXbar_portsDIO_filtered_1_valid ; 
  assign  tlMasterXbar_in_1_d_bits_opcode = tlMasterXbar_portsDIO_filtered_1_bits_opcode ; 
  assign  tlMasterXbar_in_1_d_bits_param = tlMasterXbar_portsDIO_filtered_1_bits_param ; 
  assign  tlMasterXbar_in_1_d_bits_size = tlMasterXbar_portsDIO_filtered_1_bits_size ; 
    wire tlMasterXbar_in_1_d_bits_source = tlMasterXbar_portsDIO_filtered_1_bits_source ; 
  assign  tlMasterXbar_in_1_d_bits_sink = tlMasterXbar_portsDIO_filtered_1_bits_sink ; 
  assign  tlMasterXbar_in_1_d_bits_denied = tlMasterXbar_portsDIO_filtered_1_bits_denied ; 
  assign  tlMasterXbar_in_1_d_bits_data = tlMasterXbar_portsDIO_filtered_1_bits_data ; 
  assign  tlMasterXbar_in_1_d_bits_corrupt = tlMasterXbar_portsDIO_filtered_1_bits_corrupt ; 
  assign  tlMasterXbar_portsDIO_filtered_0_valid = tlMasterXbar_out_0_d_valid & tlMasterXbar_requestDOI_0_0 ; 
  assign  tlMasterXbar_portsDIO_filtered_1_valid = tlMasterXbar_out_0_d_valid & tlMasterXbar_requestDOI_0_1 ; 
  assign  tlMasterXbar_out_0_d_ready = tlMasterXbar_requestDOI_0_0 & tlMasterXbar_portsDIO_filtered_0_ready | tlMasterXbar_requestDOI_0_1 ; reg[9:0] tlMasterXbar_beatsLeft ; 
    wire tlMasterXbar_idle = tlMasterXbar_beatsLeft ==10'h0; 
    wire tlMasterXbar_latch = tlMasterXbar_idle & tlMasterXbar_out_0_a_ready ; 
    wire[1:0] tlMasterXbar_readys_valid ={ tlMasterXbar_portsAOI_filtered_1_0_valid , tlMasterXbar_portsAOI_filtered_0_valid }; reg[1:0] tlMasterXbar_readys_mask ; 
    wire[3:0] tlMasterXbar_readys_filter ={ tlMasterXbar_readys_valid &~ tlMasterXbar_readys_mask , tlMasterXbar_readys_valid }; 
    wire[3:0] tlMasterXbar_readys_unready ={ tlMasterXbar_readys_mask [1], tlMasterXbar_readys_filter [3]| tlMasterXbar_readys_mask [0], tlMasterXbar_readys_filter [2:1]| tlMasterXbar_readys_filter [3:2]}; 
    wire[1:0] tlMasterXbar_readys_readys =~( tlMasterXbar_readys_unready [3:2]& tlMasterXbar_readys_unready [1:0]); 
    wire tlMasterXbar_readys_0 = tlMasterXbar_readys_readys [0]; 
    wire tlMasterXbar_readys_1 = tlMasterXbar_readys_readys [1]; 
    wire tlMasterXbar_winner_0 = tlMasterXbar_readys_0 & tlMasterXbar_portsAOI_filtered_0_valid ; 
    wire tlMasterXbar_winner_1 = tlMasterXbar_readys_1 & tlMasterXbar_portsAOI_filtered_1_0_valid ; 
    wire tlMasterXbar_prefixOR_1 = tlMasterXbar_winner_0 ; 
    wire tlMasterXbar__out_0_a_valid_T = tlMasterXbar_portsAOI_filtered_0_valid | tlMasterXbar_portsAOI_filtered_1_0_valid ; 
  always @( posedge  tlMasterXbar_clock )
         begin 
             if (~ tlMasterXbar_reset & tlMasterXbar_readys_valid != tlMasterXbar_readys_valid )
                 begin 
                     if (1)$error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_reset &~(~ tlMasterXbar_prefixOR_1 |~ tlMasterXbar_winner_1 ))
                 begin 
                     if (1)$error("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_reset &~(~ tlMasterXbar__out_0_a_valid_T | tlMasterXbar_winner_0 | tlMasterXbar_winner_1 ))
                 begin 
                     if (1)$error("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
                     if (1)$fatal;
                 end 
         end
    wire[9:0] tlMasterXbar_maskedBeats_0 = tlMasterXbar_winner_0  ?  tlMasterXbar_beatsAI_0 :10'h0; 
    wire[9:0] tlMasterXbar_initBeats = tlMasterXbar_maskedBeats_0 ; 
    reg tlMasterXbar_state_0 ; 
    reg tlMasterXbar_state_1 ; 
  assign  tlMasterXbar_muxState_0 = tlMasterXbar_idle  ?  tlMasterXbar_winner_0 : tlMasterXbar_state_0 ; 
    wire tlMasterXbar_muxState_1 = tlMasterXbar_idle  ?  tlMasterXbar_winner_1 : tlMasterXbar_state_1 ; 
  assign  tlMasterXbar_out_0_a_bits_source = tlMasterXbar_muxState_0 ; 
    wire tlMasterXbar_allowed_0 = tlMasterXbar_idle  ?  tlMasterXbar_readys_0 : tlMasterXbar_state_0 ; 
    wire tlMasterXbar_allowed_1 = tlMasterXbar_idle  ?  tlMasterXbar_readys_1 : tlMasterXbar_state_1 ; 
  assign  tlMasterXbar_portsAOI_filtered_0_ready = tlMasterXbar_out_0_a_ready & tlMasterXbar_allowed_0 ; 
  assign  tlMasterXbar_portsAOI_filtered_1_0_ready = tlMasterXbar_out_0_a_ready & tlMasterXbar_allowed_1 ; 
  assign  tlMasterXbar_out_0_a_valid = tlMasterXbar_idle  ?  tlMasterXbar__out_0_a_valid_T : tlMasterXbar_state_0 & tlMasterXbar_portsAOI_filtered_0_valid | tlMasterXbar_state_1 & tlMasterXbar_portsAOI_filtered_1_0_valid ; 
  assign  tlMasterXbar_out_0_a_bits_data = tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_data :32'h0; 
  assign  tlMasterXbar_out_0_a_bits_mask =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_mask :4'h0)|{4{ tlMasterXbar_muxState_1 }}; 
  assign  tlMasterXbar_out_0_a_bits_address =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_address :32'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_address :32'h0); 
  assign  tlMasterXbar_out_0_a_bits_size =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_size :4'h0)|( tlMasterXbar_muxState_1  ? 4'h6:4'h0); 
  assign  tlMasterXbar_out_0_a_bits_param = tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_param :3'h0; 
  assign  tlMasterXbar_out_0_a_bits_opcode =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_opcode :3'h0)|{ tlMasterXbar_muxState_1 ,2'h0}; 
    wire[1:0] tlMasterXbar__readys_mask_T = tlMasterXbar_readys_readys & tlMasterXbar_readys_valid ; 
  always @( posedge  tlMasterXbar_clock )
         begin 
             if ( tlMasterXbar_reset )
                 begin  
                     tlMasterXbar_beatsLeft  <=10'h0; 
                     tlMasterXbar_readys_mask  <=2'h3; 
                     tlMasterXbar_state_0  <=1'h0; 
                     tlMasterXbar_state_1  <=1'h0;
                 end 
              else 
                 begin 
                     if ( tlMasterXbar_latch ) 
                         tlMasterXbar_beatsLeft  <= tlMasterXbar_initBeats ;
                      else  
                         tlMasterXbar_beatsLeft  <= tlMasterXbar_beatsLeft -{9'h0, tlMasterXbar_out_0_a_ready & tlMasterXbar_out_0_a_valid };
                     if ( tlMasterXbar_latch &(| tlMasterXbar_readys_valid )) 
                         tlMasterXbar_readys_mask  <= tlMasterXbar__readys_mask_T |{ tlMasterXbar__readys_mask_T [0],1'h0}; 
                     tlMasterXbar_state_0  <= tlMasterXbar_muxState_0 ; 
                     tlMasterXbar_state_1  <= tlMasterXbar_muxState_1 ;
                 end 
         end
    wire tlMasterXbar_monitor_clock;
    wire tlMasterXbar_monitor_reset;
    wire tlMasterXbar_monitor_io_in_a_ready;
    wire tlMasterXbar_monitor_io_in_a_valid;
    wire[2:0] tlMasterXbar_monitor_io_in_a_bits_opcode;
    wire[2:0] tlMasterXbar_monitor_io_in_a_bits_param;
    wire[3:0] tlMasterXbar_monitor_io_in_a_bits_size;
    wire[31:0] tlMasterXbar_monitor_io_in_a_bits_address;
    wire[3:0] tlMasterXbar_monitor_io_in_a_bits_mask;
    wire tlMasterXbar_monitor_io_in_d_ready;
    wire tlMasterXbar_monitor_io_in_d_valid;
    wire[2:0] tlMasterXbar_monitor_io_in_d_bits_opcode;
    wire[1:0] tlMasterXbar_monitor_io_in_d_bits_param;
    wire[3:0] tlMasterXbar_monitor_io_in_d_bits_size;
    wire tlMasterXbar_monitor_io_in_d_bits_sink;
    wire tlMasterXbar_monitor_io_in_d_bits_denied;
    wire tlMasterXbar_monitor_io_in_d_bits_corrupt;

    wire[31:0] tlMasterXbar_monitor__plusarg_reader_1_out ; 
    wire[31:0] tlMasterXbar_monitor__plusarg_reader_out ; 
    wire tlMasterXbar_monitor_c_first =1'h1; 
    wire tlMasterXbar_monitor_c_first_last =1'h1; 
    wire tlMasterXbar_monitor_sink_ok =1'h0; 
    wire tlMasterXbar_monitor_c_first_beats1_opdata =1'h0; 
    wire tlMasterXbar_monitor_c_first_done =1'h0; 
    wire tlMasterXbar_monitor_c_set =1'h0; 
    wire tlMasterXbar_monitor_c_set_wo_ready =1'h0; 
    wire tlMasterXbar_monitor_c_probe_ack =1'h0; 
    wire tlMasterXbar_monitor_same_cycle_resp_1 =1'h0; 
    wire[9:0] tlMasterXbar_monitor_c_first_counter1 =10'h3FF; 
    wire[2:0] tlMasterXbar_monitor_responseMap_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMap_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMap_5 =3'h2; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_5 =3'h2; 
    wire[2:0] tlMasterXbar_monitor_responseMap_6 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_responseMap_7 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_7 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_6 =3'h5; 
    wire[3:0] tlMasterXbar_monitor_c_opcodes_set =4'h0; 
    wire[3:0] tlMasterXbar_monitor_c_opcodes_set_interm =4'h0; 
    wire[7:0] tlMasterXbar_monitor_c_sizes_set =8'h0; 
    wire[9:0] tlMasterXbar_monitor_c_first_beats1_decode =10'h0; 
    wire[9:0] tlMasterXbar_monitor_c_first_beats1 =10'h0; 
    wire[9:0] tlMasterXbar_monitor_c_first_count =10'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMap_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMap_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMap_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_4 =3'h1; 
    wire[4:0] tlMasterXbar_monitor_c_sizes_set_interm =5'h0; 
    wire[26:0] tlMasterXbar_monitor__GEN ={23'h0, tlMasterXbar_monitor_io_in_a_bits_size }; 
    wire[26:0] tlMasterXbar_monitor__is_aligned_mask_T_1 =27'hFFF<< tlMasterXbar_monitor__GEN ; 
    wire[11:0] tlMasterXbar_monitor_is_aligned_mask =~( tlMasterXbar_monitor__is_aligned_mask_T_1 [11:0]); 
    wire tlMasterXbar_monitor_is_aligned =( tlMasterXbar_monitor_io_in_a_bits_address [11:0]& tlMasterXbar_monitor_is_aligned_mask )==12'h0; 
    wire tlMasterXbar_monitor_mask_sizeOH_shiftAmount = tlMasterXbar_monitor_io_in_a_bits_size [0]; 
    wire[1:0] tlMasterXbar_monitor_mask_sizeOH ={ tlMasterXbar_monitor_mask_sizeOH_shiftAmount ,1'h1}; 
    wire tlMasterXbar_monitor_mask_size = tlMasterXbar_monitor_mask_sizeOH [1]; 
    wire tlMasterXbar_monitor_mask_bit = tlMasterXbar_monitor_io_in_a_bits_address [1]; 
    wire tlMasterXbar_monitor_mask_eq_1 = tlMasterXbar_monitor_mask_bit ; 
    wire tlMasterXbar_monitor_mask_nbit =~ tlMasterXbar_monitor_mask_bit ; 
    wire tlMasterXbar_monitor_mask_eq = tlMasterXbar_monitor_mask_nbit ; 
    wire tlMasterXbar_monitor_mask_acc =(|( tlMasterXbar_monitor_io_in_a_bits_size [3:1]))| tlMasterXbar_monitor_mask_size & tlMasterXbar_monitor_mask_eq ; 
    wire tlMasterXbar_monitor_mask_acc_1 =(|( tlMasterXbar_monitor_io_in_a_bits_size [3:1]))| tlMasterXbar_monitor_mask_size & tlMasterXbar_monitor_mask_eq_1 ; 
    wire tlMasterXbar_monitor_mask_size_1 = tlMasterXbar_monitor_mask_sizeOH [0]; 
    wire tlMasterXbar_monitor_mask_bit_1 = tlMasterXbar_monitor_io_in_a_bits_address [0]; 
    wire tlMasterXbar_monitor_mask_nbit_1 =~ tlMasterXbar_monitor_mask_bit_1 ; 
    wire tlMasterXbar_monitor_mask_eq_2 = tlMasterXbar_monitor_mask_eq & tlMasterXbar_monitor_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_2 = tlMasterXbar_monitor_mask_acc | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_2 ; 
    wire tlMasterXbar_monitor_mask_eq_3 = tlMasterXbar_monitor_mask_eq & tlMasterXbar_monitor_mask_bit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_3 = tlMasterXbar_monitor_mask_acc | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_3 ; 
    wire tlMasterXbar_monitor_mask_eq_4 = tlMasterXbar_monitor_mask_eq_1 & tlMasterXbar_monitor_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_4 = tlMasterXbar_monitor_mask_acc_1 | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_4 ; 
    wire tlMasterXbar_monitor_mask_eq_5 = tlMasterXbar_monitor_mask_eq_1 & tlMasterXbar_monitor_mask_bit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_5 = tlMasterXbar_monitor_mask_acc_1 | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_5 ; 
    wire[1:0] tlMasterXbar_monitor_mask_lo ={ tlMasterXbar_monitor_mask_acc_3 , tlMasterXbar_monitor_mask_acc_2 }; 
    wire[1:0] tlMasterXbar_monitor_mask_hi ={ tlMasterXbar_monitor_mask_acc_5 , tlMasterXbar_monitor_mask_acc_4 }; 
    wire[3:0] tlMasterXbar_monitor_mask ={ tlMasterXbar_monitor_mask_hi , tlMasterXbar_monitor_mask_lo }; 
    wire tlMasterXbar_monitor__GEN_0 = tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor_d_release_ack ; 
  assign  tlMasterXbar_monitor_d_release_ack = tlMasterXbar_monitor__GEN_0 ; 
    wire tlMasterXbar_monitor_d_release_ack_1 ; 
  assign  tlMasterXbar_monitor_d_release_ack_1 = tlMasterXbar_monitor__GEN_0 ; 
    wire tlMasterXbar_monitor__a_first_T_1 = tlMasterXbar_monitor_io_in_a_ready & tlMasterXbar_monitor_io_in_a_valid ; 
    wire[26:0] tlMasterXbar_monitor__a_first_beats1_decode_T_1 =27'hFFF<< tlMasterXbar_monitor__GEN ; 
    wire[9:0] tlMasterXbar_monitor_a_first_beats1_decode =~( tlMasterXbar_monitor__a_first_beats1_decode_T_1 [11:2]); 
    wire tlMasterXbar_monitor_a_first_beats1_opdata =~( tlMasterXbar_monitor_io_in_a_bits_opcode [2]); 
    wire[9:0] tlMasterXbar_monitor_a_first_beats1 = tlMasterXbar_monitor_a_first_beats1_opdata  ?  tlMasterXbar_monitor_a_first_beats1_decode :10'h0; reg[9:0] tlMasterXbar_monitor_a_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_a_first_counter1 = tlMasterXbar_monitor_a_first_counter -10'h1; 
    wire tlMasterXbar_monitor_a_first = tlMasterXbar_monitor_a_first_counter ==10'h0; 
    wire tlMasterXbar_monitor_a_first_last = tlMasterXbar_monitor_a_first_counter ==10'h1| tlMasterXbar_monitor_a_first_beats1 ==10'h0; 
    wire tlMasterXbar_monitor_a_first_done = tlMasterXbar_monitor_a_first_last & tlMasterXbar_monitor__a_first_T_1 ; 
    wire[9:0] tlMasterXbar_monitor_a_first_count = tlMasterXbar_monitor_a_first_beats1 &~ tlMasterXbar_monitor_a_first_counter1 ; reg[2:0] tlMasterXbar_monitor_opcode ; reg[2:0] tlMasterXbar_monitor_param ; reg[3:0] tlMasterXbar_monitor_size ; reg[31:0] tlMasterXbar_monitor_address ; 
    wire tlMasterXbar_monitor__d_first_T_2 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_1 ={23'h0, tlMasterXbar_monitor_io_in_d_bits_size }; 
    wire[26:0] tlMasterXbar_monitor__d_first_beats1_decode_T_1 =27'hFFF<< tlMasterXbar_monitor__GEN_1 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_beats1_decode =~( tlMasterXbar_monitor__d_first_beats1_decode_T_1 [11:2]); 
    wire tlMasterXbar_monitor_d_first_beats1_opdata = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire tlMasterXbar_monitor_d_first_beats1_opdata_1 = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire tlMasterXbar_monitor_d_first_beats1_opdata_2 = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire[9:0] tlMasterXbar_monitor_d_first_beats1 = tlMasterXbar_monitor_d_first_beats1_opdata  ?  tlMasterXbar_monitor_d_first_beats1_decode :10'h0; reg[9:0] tlMasterXbar_monitor_d_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_d_first_counter1 = tlMasterXbar_monitor_d_first_counter -10'h1; 
    wire tlMasterXbar_monitor_d_first = tlMasterXbar_monitor_d_first_counter ==10'h0; 
    wire tlMasterXbar_monitor_d_first_last = tlMasterXbar_monitor_d_first_counter ==10'h1| tlMasterXbar_monitor_d_first_beats1 ==10'h0; 
    wire tlMasterXbar_monitor_d_first_done = tlMasterXbar_monitor_d_first_last & tlMasterXbar_monitor__d_first_T_2 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_count = tlMasterXbar_monitor_d_first_beats1 &~ tlMasterXbar_monitor_d_first_counter1 ; reg[2:0] tlMasterXbar_monitor_opcode_1 ; reg[1:0] tlMasterXbar_monitor_param_1 ; reg[3:0] tlMasterXbar_monitor_size_1 ; 
    reg tlMasterXbar_monitor_sink ; 
    reg tlMasterXbar_monitor_denied ; 
    reg tlMasterXbar_monitor_inflight ; reg[3:0] tlMasterXbar_monitor_inflight_opcodes ; reg[7:0] tlMasterXbar_monitor_inflight_sizes ; 
    wire[26:0] tlMasterXbar_monitor__a_first_beats1_decode_T_5 =27'hFFF<< tlMasterXbar_monitor__GEN ; 
    wire[9:0] tlMasterXbar_monitor_a_first_beats1_decode_1 =~( tlMasterXbar_monitor__a_first_beats1_decode_T_5 [11:2]); 
    wire tlMasterXbar_monitor_a_first_beats1_opdata_1 =~( tlMasterXbar_monitor_io_in_a_bits_opcode [2]); 
    wire[9:0] tlMasterXbar_monitor_a_first_beats1_1 = tlMasterXbar_monitor_a_first_beats1_opdata_1  ?  tlMasterXbar_monitor_a_first_beats1_decode_1 :10'h0; reg[9:0] tlMasterXbar_monitor_a_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor_a_first_counter1_1 = tlMasterXbar_monitor_a_first_counter_1 -10'h1; 
    wire tlMasterXbar_monitor_a_first_1 = tlMasterXbar_monitor_a_first_counter_1 ==10'h0; 
    wire tlMasterXbar_monitor_a_first_last_1 = tlMasterXbar_monitor_a_first_counter_1 ==10'h1| tlMasterXbar_monitor_a_first_beats1_1 ==10'h0; 
    wire tlMasterXbar_monitor_a_first_done_1 = tlMasterXbar_monitor_a_first_last_1 & tlMasterXbar_monitor__a_first_T_1 ; 
    wire[9:0] tlMasterXbar_monitor_a_first_count_1 = tlMasterXbar_monitor_a_first_beats1_1 &~ tlMasterXbar_monitor_a_first_counter1_1 ; 
    wire[26:0] tlMasterXbar_monitor__d_first_beats1_decode_T_5 =27'hFFF<< tlMasterXbar_monitor__GEN_1 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_beats1_decode_1 =~( tlMasterXbar_monitor__d_first_beats1_decode_T_5 [11:2]); 
    wire[9:0] tlMasterXbar_monitor_d_first_beats1_1 = tlMasterXbar_monitor_d_first_beats1_opdata_1  ?  tlMasterXbar_monitor_d_first_beats1_decode_1 :10'h0; reg[9:0] tlMasterXbar_monitor_d_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_counter1_1 = tlMasterXbar_monitor_d_first_counter_1 -10'h1; 
    wire tlMasterXbar_monitor_d_first_1 = tlMasterXbar_monitor_d_first_counter_1 ==10'h0; 
    wire tlMasterXbar_monitor_d_first_last_1 = tlMasterXbar_monitor_d_first_counter_1 ==10'h1| tlMasterXbar_monitor_d_first_beats1_1 ==10'h0; 
    wire tlMasterXbar_monitor_d_first_done_1 = tlMasterXbar_monitor_d_first_last_1 & tlMasterXbar_monitor__d_first_T_2 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_count_1 = tlMasterXbar_monitor_d_first_beats1_1 &~ tlMasterXbar_monitor_d_first_counter1_1 ; 
    wire[3:0] tlMasterXbar_monitor_a_opcode_lookup ={1'h0, tlMasterXbar_monitor_inflight_opcodes [3:1]}; 
    wire[7:0] tlMasterXbar_monitor_a_size_lookup ={1'h0, tlMasterXbar_monitor_inflight_sizes [7:1]}; 
    wire tlMasterXbar_monitor__same_cycle_resp_T_1 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_a_first_1 ; 
    wire tlMasterXbar_monitor_a_set_wo_ready ; 
  assign  tlMasterXbar_monitor_a_set_wo_ready = tlMasterXbar_monitor__same_cycle_resp_T_1 ; 
    wire tlMasterXbar_monitor_same_cycle_resp ; 
  assign  tlMasterXbar_monitor_same_cycle_resp = tlMasterXbar_monitor__same_cycle_resp_T_1 ; 
    wire tlMasterXbar_monitor_a_set = tlMasterXbar_monitor__a_first_T_1 & tlMasterXbar_monitor_a_first_1 ; 
    wire[3:0] tlMasterXbar_monitor_a_opcodes_set_interm = tlMasterXbar_monitor_a_set  ? { tlMasterXbar_monitor_io_in_a_bits_opcode ,1'h1}:4'h0; 
    wire[4:0] tlMasterXbar_monitor_a_sizes_set_interm = tlMasterXbar_monitor_a_set  ? { tlMasterXbar_monitor_io_in_a_bits_size ,1'h1}:5'h0; 
    wire[3:0] tlMasterXbar_monitor_a_opcodes_set = tlMasterXbar_monitor_a_set  ?  tlMasterXbar_monitor_a_opcodes_set_interm :4'h0; 
    wire[7:0] tlMasterXbar_monitor_a_sizes_set = tlMasterXbar_monitor_a_set  ? {3'h0, tlMasterXbar_monitor_a_sizes_set_interm }:8'h0; 
    wire tlMasterXbar_monitor__GEN_2 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_1 ; 
    wire tlMasterXbar_monitor_d_clr_wo_ready = tlMasterXbar_monitor__GEN_2 &~ tlMasterXbar_monitor_d_release_ack ; 
    wire tlMasterXbar_monitor_d_clr = tlMasterXbar_monitor__d_first_T_2 & tlMasterXbar_monitor_d_first_1 &~ tlMasterXbar_monitor_d_release_ack ; 
    wire[3:0] tlMasterXbar_monitor_d_opcodes_clr ={4{ tlMasterXbar_monitor_d_clr }}; 
    wire[7:0] tlMasterXbar_monitor_d_sizes_clr ={8{ tlMasterXbar_monitor_d_clr }}; reg[2:0] tlMasterXbar_monitor_casez_tmp ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_io_in_a_bits_opcode )
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp  =3'h0;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp  =3'h0;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp  =3'h1;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp  =3'h1;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp  =3'h1;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp  =3'h2;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp  =3'h4;
              default : 
                  tlMasterXbar_monitor_casez_tmp  =3'h4;endcase
         end
  reg[2:0] tlMasterXbar_monitor_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_io_in_a_bits_opcode )
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h0;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h0;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h1;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h1;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h1;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h2;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h5;
              default : 
                  tlMasterXbar_monitor_casez_tmp_0  =3'h4;endcase
         end
  reg[2:0] tlMasterXbar_monitor_casez_tmp_1 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h0;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h0;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h1;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h1;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h1;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h2;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h4;
              default : 
                  tlMasterXbar_monitor_casez_tmp_1  =3'h4;endcase
         end
  reg[2:0] tlMasterXbar_monitor_casez_tmp_2 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h0;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h0;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h1;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h1;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h1;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h2;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h5;
              default : 
                  tlMasterXbar_monitor_casez_tmp_2  =3'h4;endcase
         end
  reg[31:0] tlMasterXbar_monitor_watchdog ; 
    reg tlMasterXbar_monitor_inflight_1 ; reg[3:0] tlMasterXbar_monitor_inflight_opcodes_1 ; reg[7:0] tlMasterXbar_monitor_inflight_sizes_1 ; 
    wire[26:0] tlMasterXbar_monitor__d_first_beats1_decode_T_9 =27'hFFF<< tlMasterXbar_monitor__GEN_1 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_beats1_decode_2 =~( tlMasterXbar_monitor__d_first_beats1_decode_T_9 [11:2]); 
    wire[9:0] tlMasterXbar_monitor_d_first_beats1_2 = tlMasterXbar_monitor_d_first_beats1_opdata_2  ?  tlMasterXbar_monitor_d_first_beats1_decode_2 :10'h0; reg[9:0] tlMasterXbar_monitor_d_first_counter_2 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_counter1_2 = tlMasterXbar_monitor_d_first_counter_2 -10'h1; 
    wire tlMasterXbar_monitor_d_first_2 = tlMasterXbar_monitor_d_first_counter_2 ==10'h0; 
    wire tlMasterXbar_monitor_d_first_last_2 = tlMasterXbar_monitor_d_first_counter_2 ==10'h1| tlMasterXbar_monitor_d_first_beats1_2 ==10'h0; 
    wire tlMasterXbar_monitor_d_first_done_2 = tlMasterXbar_monitor_d_first_last_2 & tlMasterXbar_monitor__d_first_T_2 ; 
    wire[9:0] tlMasterXbar_monitor_d_first_count_2 = tlMasterXbar_monitor_d_first_beats1_2 &~ tlMasterXbar_monitor_d_first_counter1_2 ; 
    wire[3:0] tlMasterXbar_monitor_c_opcode_lookup ={1'h0, tlMasterXbar_monitor_inflight_opcodes_1 [3:1]}; 
    wire[7:0] tlMasterXbar_monitor_c_size_lookup ={1'h0, tlMasterXbar_monitor_inflight_sizes_1 [7:1]}; 
    wire tlMasterXbar_monitor_d_clr_wo_ready_1 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_2 & tlMasterXbar_monitor_d_release_ack_1 ; 
    wire tlMasterXbar_monitor_d_clr_1 = tlMasterXbar_monitor__d_first_T_2 & tlMasterXbar_monitor_d_first_2 & tlMasterXbar_monitor_d_release_ack_1 ; 
    wire[3:0] tlMasterXbar_monitor_d_opcodes_clr_1 ={4{ tlMasterXbar_monitor_d_clr_1 }}; 
    wire[7:0] tlMasterXbar_monitor_d_sizes_clr_1 ={8{ tlMasterXbar_monitor_d_clr_1 }}; reg[31:0] tlMasterXbar_monitor_watchdog_1 ; 
    wire tlMasterXbar_monitor__GEN_3 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h6&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_4 = tlMasterXbar_monitor_io_in_a_bits_param >3'h2; 
    wire tlMasterXbar_monitor__GEN_5 = tlMasterXbar_monitor_io_in_a_bits_mask !=4'hF; 
    wire tlMasterXbar_monitor__GEN_6 = tlMasterXbar_monitor_io_in_a_valid &(& tlMasterXbar_monitor_io_in_a_bits_opcode )&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_7 = tlMasterXbar_monitor_io_in_a_bits_size <4'hD; 
    wire tlMasterXbar_monitor__GEN_8 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h4&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_9 ={ tlMasterXbar_monitor_io_in_a_bits_address [31:14],~( tlMasterXbar_monitor_io_in_a_bits_address [13:12])}==20'h0; 
    wire tlMasterXbar_monitor__GEN_10 = tlMasterXbar_monitor__GEN_7 & tlMasterXbar_monitor__GEN_9 ; 
    wire tlMasterXbar_monitor__GEN_11 = tlMasterXbar_monitor_io_in_a_bits_size <4'h7; 
    wire tlMasterXbar_monitor__GEN_12 = tlMasterXbar_monitor_io_in_a_bits_address [31:12]==20'h0; 
    wire tlMasterXbar_monitor__GEN_13 ={ tlMasterXbar_monitor_io_in_a_bits_address [31:26], tlMasterXbar_monitor_io_in_a_bits_address [25:16]^10'h200}==16'h0; 
    wire tlMasterXbar_monitor__GEN_14 ={ tlMasterXbar_monitor_io_in_a_bits_address [31:28],~( tlMasterXbar_monitor_io_in_a_bits_address [27:26])}==6'h0; 
    wire tlMasterXbar_monitor__GEN_15 ={ tlMasterXbar_monitor_io_in_a_bits_address [31],~( tlMasterXbar_monitor_io_in_a_bits_address [30:29])}==3'h0; 
    wire tlMasterXbar_monitor__GEN_16 = tlMasterXbar_monitor_io_in_a_bits_address [31:14]==18'h20000; 
    wire tlMasterXbar_monitor__GEN_17 = tlMasterXbar_monitor_io_in_a_bits_mask != tlMasterXbar_monitor_mask ; 
    wire tlMasterXbar_monitor__GEN_18 = tlMasterXbar_monitor__GEN_7 &( tlMasterXbar_monitor__GEN_10 | tlMasterXbar_monitor__GEN_11 &( tlMasterXbar_monitor__GEN_12 | tlMasterXbar_monitor__GEN_13 | tlMasterXbar_monitor__GEN_14 | tlMasterXbar_monitor__GEN_16 )| tlMasterXbar_monitor_io_in_a_bits_size <4'h9& tlMasterXbar_monitor__GEN_15 ); 
    wire tlMasterXbar_monitor__GEN_19 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h0&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_20 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h1&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_21 = tlMasterXbar_monitor__GEN_7 & tlMasterXbar_monitor_io_in_a_bits_size <4'h3&( tlMasterXbar_monitor__GEN_12 | tlMasterXbar_monitor__GEN_9 | tlMasterXbar_monitor__GEN_13 | tlMasterXbar_monitor__GEN_14 | tlMasterXbar_monitor__GEN_16 ); 
    wire tlMasterXbar_monitor__GEN_22 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h2&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_23 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h3&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_24 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h5&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_25 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor__GEN_0 &~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_26 = tlMasterXbar_monitor_io_in_d_bits_size [3:1]==3'h0; 
    wire tlMasterXbar_monitor__GEN_27 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h4&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_28 = tlMasterXbar_monitor_io_in_d_bits_param ==2'h2; 
    wire tlMasterXbar_monitor__GEN_29 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h5&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_30 =~ tlMasterXbar_monitor_io_in_d_bits_denied | tlMasterXbar_monitor_io_in_d_bits_corrupt ; 
    wire tlMasterXbar_monitor__GEN_31 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h0&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_32 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h1&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_33 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h2&~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_34 = tlMasterXbar_monitor_io_in_a_valid &~ tlMasterXbar_monitor_a_first &~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_35 = tlMasterXbar_monitor_io_in_d_valid &~ tlMasterXbar_monitor_d_first &~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_36 = tlMasterXbar_monitor_d_clr_wo_ready & tlMasterXbar_monitor_same_cycle_resp &~ tlMasterXbar_monitor_reset ; 
    wire tlMasterXbar_monitor__GEN_37 = tlMasterXbar_monitor_d_clr_wo_ready &~ tlMasterXbar_monitor_same_cycle_resp &~ tlMasterXbar_monitor_reset ; 
    wire[7:0] tlMasterXbar_monitor__GEN_38 ={4'h0, tlMasterXbar_monitor_io_in_d_bits_size }; 
    wire tlMasterXbar_monitor__GEN_39 = tlMasterXbar_monitor_d_clr_wo_ready_1 &~ tlMasterXbar_monitor_reset ; 
  always @( posedge  tlMasterXbar_monitor_clock )
         begin 
             if ( tlMasterXbar_monitor__GEN_3 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                     if (1)$error("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 &~(|( tlMasterXbar_monitor_io_in_a_bits_size [3:1])))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor__GEN_4 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor__GEN_5 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_6 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                     if (1)$error("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_6 &~(|( tlMasterXbar_monitor_io_in_a_bits_size [3:1])))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_6 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_6 & tlMasterXbar_monitor__GEN_4 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_6 &~(| tlMasterXbar_monitor_io_in_a_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_6 & tlMasterXbar_monitor__GEN_5 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_8 &~ tlMasterXbar_monitor__GEN_7 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_8 &~( tlMasterXbar_monitor__GEN_10 | tlMasterXbar_monitor__GEN_11 &( tlMasterXbar_monitor__GEN_12 |{ tlMasterXbar_monitor_io_in_a_bits_address [31:17],~( tlMasterXbar_monitor_io_in_a_bits_address [16])}==16'h0| tlMasterXbar_monitor__GEN_13 | tlMasterXbar_monitor__GEN_14 | tlMasterXbar_monitor__GEN_15 | tlMasterXbar_monitor__GEN_16 )))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_8 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_8 &(| tlMasterXbar_monitor_io_in_a_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_8 & tlMasterXbar_monitor__GEN_17 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_19 &~ tlMasterXbar_monitor__GEN_18 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_19 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_19 &(| tlMasterXbar_monitor_io_in_a_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_19 & tlMasterXbar_monitor__GEN_17 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_20 &~ tlMasterXbar_monitor__GEN_18 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_20 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_20 &(| tlMasterXbar_monitor_io_in_a_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_20 &(|( tlMasterXbar_monitor_io_in_a_bits_mask &~ tlMasterXbar_monitor_mask )))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_22 &~ tlMasterXbar_monitor__GEN_21 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_22 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_22 & tlMasterXbar_monitor_io_in_a_bits_param >3'h4)
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_22 & tlMasterXbar_monitor__GEN_17 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_23 &~ tlMasterXbar_monitor__GEN_21 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_23 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_23 & tlMasterXbar_monitor_io_in_a_bits_param [2])
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_23 & tlMasterXbar_monitor__GEN_17 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_24 &~( tlMasterXbar_monitor__GEN_7 & tlMasterXbar_monitor__GEN_10 ))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_24 &~ tlMasterXbar_monitor_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_24 &(|( tlMasterXbar_monitor_io_in_a_bits_param [2:1])))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_24 & tlMasterXbar_monitor__GEN_17 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_d_valid &~ tlMasterXbar_monitor_reset &(& tlMasterXbar_monitor_io_in_d_bits_opcode ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_25 & tlMasterXbar_monitor__GEN_26 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_25 &(| tlMasterXbar_monitor_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_25 & tlMasterXbar_monitor_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_25 & tlMasterXbar_monitor_io_in_d_bits_denied )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_27 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_27 & tlMasterXbar_monitor__GEN_26 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_27 &(& tlMasterXbar_monitor_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_27 & tlMasterXbar_monitor__GEN_28 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_27 & tlMasterXbar_monitor_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_29 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_29 & tlMasterXbar_monitor__GEN_26 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_29 &(& tlMasterXbar_monitor_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_29 & tlMasterXbar_monitor__GEN_28 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_29 &~ tlMasterXbar_monitor__GEN_30 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_31 &(| tlMasterXbar_monitor_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_31 & tlMasterXbar_monitor_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_32 &(| tlMasterXbar_monitor_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_32 &~ tlMasterXbar_monitor__GEN_30 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_33 &(| tlMasterXbar_monitor_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_33 & tlMasterXbar_monitor_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_34 & tlMasterXbar_monitor_io_in_a_bits_opcode != tlMasterXbar_monitor_opcode )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_34 & tlMasterXbar_monitor_io_in_a_bits_param != tlMasterXbar_monitor_param )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_34 & tlMasterXbar_monitor_io_in_a_bits_size != tlMasterXbar_monitor_size )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_34 & tlMasterXbar_monitor_io_in_a_bits_address != tlMasterXbar_monitor_address )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_35 & tlMasterXbar_monitor_io_in_d_bits_opcode != tlMasterXbar_monitor_opcode_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_35 & tlMasterXbar_monitor_io_in_d_bits_param != tlMasterXbar_monitor_param_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_35 & tlMasterXbar_monitor_io_in_d_bits_size != tlMasterXbar_monitor_size_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_35 & tlMasterXbar_monitor_io_in_d_bits_sink != tlMasterXbar_monitor_sink )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_35 & tlMasterXbar_monitor_io_in_d_bits_denied != tlMasterXbar_monitor_denied )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_a_set &~ tlMasterXbar_monitor_reset & tlMasterXbar_monitor_inflight )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_d_clr_wo_ready &~ tlMasterXbar_monitor_reset &~( tlMasterXbar_monitor_inflight | tlMasterXbar_monitor_same_cycle_resp ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 &~( tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp | tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp_0 ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 & tlMasterXbar_monitor_io_in_a_bits_size != tlMasterXbar_monitor_io_in_d_bits_size )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_37 &~( tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp_1 | tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp_2 ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_37 & tlMasterXbar_monitor__GEN_38 != tlMasterXbar_monitor_a_size_lookup )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_2 & tlMasterXbar_monitor_a_first_1 & tlMasterXbar_monitor_io_in_a_valid &~ tlMasterXbar_monitor_d_release_ack &~ tlMasterXbar_monitor_reset &~(~ tlMasterXbar_monitor_io_in_d_ready | tlMasterXbar_monitor_io_in_a_ready ))
                 begin 
                     if (1)$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_monitor_reset &~( tlMasterXbar_monitor_a_set_wo_ready != tlMasterXbar_monitor_d_clr_wo_ready |~ tlMasterXbar_monitor_a_set_wo_ready ))
                 begin 
                     if (1)$error("Assertion failed: 'A' and 'D' concurrent, despite minlatency 4 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_monitor_reset &~(~ tlMasterXbar_monitor_inflight | tlMasterXbar_monitor__plusarg_reader_out ==32'h0| tlMasterXbar_monitor_watchdog < tlMasterXbar_monitor__plusarg_reader_out ))
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_39 &~ tlMasterXbar_monitor_inflight_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_39 & tlMasterXbar_monitor__GEN_38 != tlMasterXbar_monitor_c_size_lookup )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_monitor_reset &~(~ tlMasterXbar_monitor_inflight_1 | tlMasterXbar_monitor__plusarg_reader_1_out ==32'h0| tlMasterXbar_monitor_watchdog_1 < tlMasterXbar_monitor__plusarg_reader_1_out ))
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
         end
  always @( posedge  tlMasterXbar_monitor_clock )
         begin 
             if ( tlMasterXbar_monitor_reset )
                 begin  
                     tlMasterXbar_monitor_a_first_counter  <=10'h0; 
                     tlMasterXbar_monitor_d_first_counter  <=10'h0; 
                     tlMasterXbar_monitor_inflight  <=1'h0; 
                     tlMasterXbar_monitor_inflight_opcodes  <=4'h0; 
                     tlMasterXbar_monitor_inflight_sizes  <=8'h0; 
                     tlMasterXbar_monitor_a_first_counter_1  <=10'h0; 
                     tlMasterXbar_monitor_d_first_counter_1  <=10'h0; 
                     tlMasterXbar_monitor_watchdog  <=32'h0; 
                     tlMasterXbar_monitor_inflight_1  <=1'h0; 
                     tlMasterXbar_monitor_inflight_opcodes_1  <=4'h0; 
                     tlMasterXbar_monitor_inflight_sizes_1  <=8'h0; 
                     tlMasterXbar_monitor_d_first_counter_2  <=10'h0; 
                     tlMasterXbar_monitor_watchdog_1  <=32'h0;
                 end 
              else 
                 begin 
                     if ( tlMasterXbar_monitor__a_first_T_1 )
                         begin 
                             if ( tlMasterXbar_monitor_a_first ) 
                                 tlMasterXbar_monitor_a_first_counter  <= tlMasterXbar_monitor_a_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_a_first_counter  <= tlMasterXbar_monitor_a_first_counter1 ;
                             if ( tlMasterXbar_monitor_a_first_1 ) 
                                 tlMasterXbar_monitor_a_first_counter_1  <= tlMasterXbar_monitor_a_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_a_first_counter_1  <= tlMasterXbar_monitor_a_first_counter1_1 ;
                         end 
                     if ( tlMasterXbar_monitor__d_first_T_2 )
                         begin 
                             if ( tlMasterXbar_monitor_d_first ) 
                                 tlMasterXbar_monitor_d_first_counter  <= tlMasterXbar_monitor_d_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter  <= tlMasterXbar_monitor_d_first_counter1 ;
                             if ( tlMasterXbar_monitor_d_first_1 ) 
                                 tlMasterXbar_monitor_d_first_counter_1  <= tlMasterXbar_monitor_d_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter_1  <= tlMasterXbar_monitor_d_first_counter1_1 ;
                             if ( tlMasterXbar_monitor_d_first_2 ) 
                                 tlMasterXbar_monitor_d_first_counter_2  <= tlMasterXbar_monitor_d_first_beats1_2 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter_2  <= tlMasterXbar_monitor_d_first_counter1_2 ; 
                             tlMasterXbar_monitor_watchdog_1  <=32'h0;
                         end 
                      else  
                         tlMasterXbar_monitor_watchdog_1  <= tlMasterXbar_monitor_watchdog_1 +32'h1; 
                     tlMasterXbar_monitor_inflight  <=( tlMasterXbar_monitor_inflight | tlMasterXbar_monitor_a_set )&~ tlMasterXbar_monitor_d_clr ; 
                     tlMasterXbar_monitor_inflight_opcodes  <=( tlMasterXbar_monitor_inflight_opcodes | tlMasterXbar_monitor_a_opcodes_set )&~ tlMasterXbar_monitor_d_opcodes_clr ; 
                     tlMasterXbar_monitor_inflight_sizes  <=( tlMasterXbar_monitor_inflight_sizes | tlMasterXbar_monitor_a_sizes_set )&~ tlMasterXbar_monitor_d_sizes_clr ;
                     if ( tlMasterXbar_monitor__a_first_T_1 | tlMasterXbar_monitor__d_first_T_2 ) 
                         tlMasterXbar_monitor_watchdog  <=32'h0;
                      else  
                         tlMasterXbar_monitor_watchdog  <= tlMasterXbar_monitor_watchdog +32'h1; 
                     tlMasterXbar_monitor_inflight_1  <= tlMasterXbar_monitor_inflight_1 &~ tlMasterXbar_monitor_d_clr_1 ; 
                     tlMasterXbar_monitor_inflight_opcodes_1  <= tlMasterXbar_monitor_inflight_opcodes_1 &~ tlMasterXbar_monitor_d_opcodes_clr_1 ; 
                     tlMasterXbar_monitor_inflight_sizes_1  <= tlMasterXbar_monitor_inflight_sizes_1 &~ tlMasterXbar_monitor_d_sizes_clr_1 ;
                 end 
             if ( tlMasterXbar_monitor__a_first_T_1 & tlMasterXbar_monitor_a_first )
                 begin  
                     tlMasterXbar_monitor_opcode  <= tlMasterXbar_monitor_io_in_a_bits_opcode ; 
                     tlMasterXbar_monitor_param  <= tlMasterXbar_monitor_io_in_a_bits_param ; 
                     tlMasterXbar_monitor_size  <= tlMasterXbar_monitor_io_in_a_bits_size ; 
                     tlMasterXbar_monitor_address  <= tlMasterXbar_monitor_io_in_a_bits_address ;
                 end 
             if ( tlMasterXbar_monitor__d_first_T_2 & tlMasterXbar_monitor_d_first )
                 begin  
                     tlMasterXbar_monitor_opcode_1  <= tlMasterXbar_monitor_io_in_d_bits_opcode ; 
                     tlMasterXbar_monitor_param_1  <= tlMasterXbar_monitor_io_in_d_bits_param ; 
                     tlMasterXbar_monitor_size_1  <= tlMasterXbar_monitor_io_in_d_bits_size ; 
                     tlMasterXbar_monitor_sink  <= tlMasterXbar_monitor_io_in_d_bits_sink ; 
                     tlMasterXbar_monitor_denied  <= tlMasterXbar_monitor_io_in_d_bits_denied ;
                 end 
         end
    plusarg_reader  #(. tlMasterXbar_monitor_DEFAULT (0),. tlMasterXbar_monitor_FORMAT ("tilelink_timeout=%d"),. tlMasterXbar_monitor_WIDTH (32)) tlMasterXbar_monitor_plusarg_reader (. out ( tlMasterXbar_monitor__plusarg_reader_out ));  
    plusarg_reader  #(. tlMasterXbar_monitor_DEFAULT (0),. tlMasterXbar_monitor_FORMAT ("tilelink_timeout=%d"),. tlMasterXbar_monitor_WIDTH (32)) tlMasterXbar_monitor_plusarg_reader_1 (. out ( tlMasterXbar_monitor__plusarg_reader_1_out ));
    assign tlMasterXbar_monitor_clock = tlMasterXbar_clock;
    assign tlMasterXbar_monitor_reset = tlMasterXbar_reset;
    assign tlMasterXbar_monitor_io_in_a_ready = tlMasterXbar_nodeIn_a_ready;
    assign tlMasterXbar_monitor_io_in_a_valid = tlMasterXbar_nodeIn_a_valid;
    assign tlMasterXbar_monitor_io_in_a_bits_opcode = tlMasterXbar_nodeIn_a_bits_opcode;
    assign tlMasterXbar_monitor_io_in_a_bits_param = tlMasterXbar_nodeIn_a_bits_param;
    assign tlMasterXbar_monitor_io_in_a_bits_size = tlMasterXbar_nodeIn_a_bits_size;
    assign tlMasterXbar_monitor_io_in_a_bits_address = tlMasterXbar_nodeIn_a_bits_address;
    assign tlMasterXbar_monitor_io_in_a_bits_mask = tlMasterXbar_nodeIn_a_bits_mask;
    assign tlMasterXbar_monitor_io_in_d_ready = tlMasterXbar_nodeIn_d_ready;
    assign tlMasterXbar_monitor_io_in_d_valid = tlMasterXbar_nodeIn_d_valid;
    assign tlMasterXbar_monitor_io_in_d_bits_opcode = tlMasterXbar_nodeIn_d_bits_opcode;
    assign tlMasterXbar_monitor_io_in_d_bits_param = tlMasterXbar_nodeIn_d_bits_param;
    assign tlMasterXbar_monitor_io_in_d_bits_size = tlMasterXbar_nodeIn_d_bits_size;
    assign tlMasterXbar_monitor_io_in_d_bits_sink = tlMasterXbar_nodeIn_d_bits_sink;
    assign tlMasterXbar_monitor_io_in_d_bits_denied = tlMasterXbar_nodeIn_d_bits_denied;
    assign tlMasterXbar_monitor_io_in_d_bits_corrupt = tlMasterXbar_nodeIn_d_bits_corrupt;
      
    wire tlMasterXbar_monitor_1_clock;
    wire tlMasterXbar_monitor_1_reset;
    wire tlMasterXbar_monitor_1_io_in_a_ready;
    wire tlMasterXbar_monitor_1_io_in_a_valid;
    wire[31:0] tlMasterXbar_monitor_1_io_in_a_bits_address;
    wire tlMasterXbar_monitor_1_io_in_d_valid;
    wire[2:0] tlMasterXbar_monitor_1_io_in_d_bits_opcode;
    wire[1:0] tlMasterXbar_monitor_1_io_in_d_bits_param;
    wire[3:0] tlMasterXbar_monitor_1_io_in_d_bits_size;
    wire tlMasterXbar_monitor_1_io_in_d_bits_sink;
    wire tlMasterXbar_monitor_1_io_in_d_bits_denied;
    wire tlMasterXbar_monitor_1_io_in_d_bits_corrupt;

    wire[31:0] tlMasterXbar_monitor_1__plusarg_reader_1_out ; 
    wire[31:0] tlMasterXbar_monitor_1__plusarg_reader_out ; 
    wire[1:0] tlMasterXbar_monitor_1_mask_lo =2'h3; 
    wire[1:0] tlMasterXbar_monitor_1_mask_hi =2'h3; 
    wire tlMasterXbar_monitor_1_mask_acc =1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc_1 =1'h1; 
    wire tlMasterXbar_monitor_1_mask_size_1 =1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc_2 =1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc_3 =1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc_4 =1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc_5 =1'h1; 
    wire tlMasterXbar_monitor_1_a_first_last =1'h1; 
    wire tlMasterXbar_monitor_1_a_first_last_1 =1'h1; 
    wire tlMasterXbar_monitor_1_c_first =1'h1; 
    wire tlMasterXbar_monitor_1_c_first_last =1'h1; 
    wire tlMasterXbar_monitor_1_mask_sizeOH_shiftAmount =1'h0; 
    wire tlMasterXbar_monitor_1_mask_size =1'h0; 
    wire tlMasterXbar_monitor_1_sink_ok =1'h0; 
    wire tlMasterXbar_monitor_1_a_first_beats1_opdata =1'h0; 
    wire tlMasterXbar_monitor_1_a_first_beats1_opdata_1 =1'h0; 
    wire tlMasterXbar_monitor_1_c_first_beats1_opdata =1'h0; 
    wire tlMasterXbar_monitor_1_c_first_done =1'h0; 
    wire tlMasterXbar_monitor_1_c_set =1'h0; 
    wire tlMasterXbar_monitor_1_c_set_wo_ready =1'h0; 
    wire tlMasterXbar_monitor_1_c_probe_ack =1'h0; 
    wire tlMasterXbar_monitor_1_same_cycle_resp_1 =1'h0; 
    wire[9:0] tlMasterXbar_monitor_1_c_first_counter1 =10'h3FF; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_6 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_7 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_7 =3'h4; 
    wire[3:0] tlMasterXbar_monitor_1_mask =4'hF; 
    wire[3:0] tlMasterXbar_monitor_1_c_opcodes_set =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1_c_opcodes_set_interm =4'h0; 
    wire[7:0] tlMasterXbar_monitor_1_c_sizes_set =8'h0; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_beats1 =10'h0; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_count =10'h0; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_beats1_1 =10'h0; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_count_1 =10'h0; 
    wire[9:0] tlMasterXbar_monitor_1_c_first_beats1_decode =10'h0; 
    wire[9:0] tlMasterXbar_monitor_1_c_first_beats1 =10'h0; 
    wire[9:0] tlMasterXbar_monitor_1_c_first_count =10'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_6 =3'h5; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_5 =3'h2; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_5 =3'h2; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_beats1_decode =10'hF; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_beats1_decode_1 =10'hF; 
    wire[1:0] tlMasterXbar_monitor_1_mask_sizeOH =2'h1; 
    wire[11:0] tlMasterXbar_monitor_1_is_aligned_mask =12'h3F; 
    wire[4:0] tlMasterXbar_monitor_1_c_sizes_set_interm =5'h0; 
    wire tlMasterXbar_monitor_1_is_aligned = tlMasterXbar_monitor_1_io_in_a_bits_address [5:0]==6'h0; 
    wire tlMasterXbar_monitor_1_mask_bit = tlMasterXbar_monitor_1_io_in_a_bits_address [1]; 
    wire tlMasterXbar_monitor_1_mask_eq_1 = tlMasterXbar_monitor_1_mask_bit ; 
    wire tlMasterXbar_monitor_1_mask_nbit =~ tlMasterXbar_monitor_1_mask_bit ; 
    wire tlMasterXbar_monitor_1_mask_eq = tlMasterXbar_monitor_1_mask_nbit ; 
    wire tlMasterXbar_monitor_1_mask_bit_1 = tlMasterXbar_monitor_1_io_in_a_bits_address [0]; 
    wire tlMasterXbar_monitor_1_mask_nbit_1 =~ tlMasterXbar_monitor_1_mask_bit_1 ; 
    wire tlMasterXbar_monitor_1_mask_eq_2 = tlMasterXbar_monitor_1_mask_eq & tlMasterXbar_monitor_1_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_1_mask_eq_3 = tlMasterXbar_monitor_1_mask_eq & tlMasterXbar_monitor_1_mask_bit_1 ; 
    wire tlMasterXbar_monitor_1_mask_eq_4 = tlMasterXbar_monitor_1_mask_eq_1 & tlMasterXbar_monitor_1_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_1_mask_eq_5 = tlMasterXbar_monitor_1_mask_eq_1 & tlMasterXbar_monitor_1_mask_bit_1 ; 
    wire tlMasterXbar_monitor_1__GEN = tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor_1_d_release_ack ; 
  assign  tlMasterXbar_monitor_1_d_release_ack = tlMasterXbar_monitor_1__GEN ; 
    wire tlMasterXbar_monitor_1_d_release_ack_1 ; 
  assign  tlMasterXbar_monitor_1_d_release_ack_1 = tlMasterXbar_monitor_1__GEN ; 
    wire tlMasterXbar_monitor_1__a_first_T_1 = tlMasterXbar_monitor_1_io_in_a_ready & tlMasterXbar_monitor_1_io_in_a_valid ; 
    wire tlMasterXbar_monitor_1_a_first_done ; 
  assign  tlMasterXbar_monitor_1_a_first_done = tlMasterXbar_monitor_1__a_first_T_1 ; 
    wire tlMasterXbar_monitor_1_a_first_done_1 ; 
  assign  tlMasterXbar_monitor_1_a_first_done_1 = tlMasterXbar_monitor_1__a_first_T_1 ; reg[9:0] tlMasterXbar_monitor_1_a_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_counter1 = tlMasterXbar_monitor_1_a_first_counter -10'h1; 
    wire tlMasterXbar_monitor_1_a_first = tlMasterXbar_monitor_1_a_first_counter ==10'h0; reg[31:0] tlMasterXbar_monitor_1_address ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_0 ={23'h0, tlMasterXbar_monitor_1_io_in_d_bits_size }; 
    wire[26:0] tlMasterXbar_monitor_1__d_first_beats1_decode_T_1 =27'hFFF<< tlMasterXbar_monitor_1__GEN_0 ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_beats1_decode =~( tlMasterXbar_monitor_1__d_first_beats1_decode_T_1 [11:2]); 
    wire tlMasterXbar_monitor_1_d_first_beats1_opdata = tlMasterXbar_monitor_1_io_in_d_bits_opcode [0]; 
    wire tlMasterXbar_monitor_1_d_first_beats1_opdata_1 = tlMasterXbar_monitor_1_io_in_d_bits_opcode [0]; 
    wire tlMasterXbar_monitor_1_d_first_beats1_opdata_2 = tlMasterXbar_monitor_1_io_in_d_bits_opcode [0]; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_beats1 = tlMasterXbar_monitor_1_d_first_beats1_opdata  ?  tlMasterXbar_monitor_1_d_first_beats1_decode :10'h0; reg[9:0] tlMasterXbar_monitor_1_d_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_counter1 = tlMasterXbar_monitor_1_d_first_counter -10'h1; 
    wire tlMasterXbar_monitor_1_d_first = tlMasterXbar_monitor_1_d_first_counter ==10'h0; 
    wire tlMasterXbar_monitor_1_d_first_last = tlMasterXbar_monitor_1_d_first_counter ==10'h1| tlMasterXbar_monitor_1_d_first_beats1 ==10'h0; 
    wire tlMasterXbar_monitor_1_d_first_done = tlMasterXbar_monitor_1_d_first_last & tlMasterXbar_monitor_1_io_in_d_valid ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_count = tlMasterXbar_monitor_1_d_first_beats1 &~ tlMasterXbar_monitor_1_d_first_counter1 ; reg[2:0] tlMasterXbar_monitor_1_opcode_1 ; reg[1:0] tlMasterXbar_monitor_1_param_1 ; reg[3:0] tlMasterXbar_monitor_1_size_1 ; 
    reg tlMasterXbar_monitor_1_sink ; 
    reg tlMasterXbar_monitor_1_denied ; 
    reg tlMasterXbar_monitor_1_inflight ; reg[3:0] tlMasterXbar_monitor_1_inflight_opcodes ; reg[7:0] tlMasterXbar_monitor_1_inflight_sizes ; reg[9:0] tlMasterXbar_monitor_1_a_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor_1_a_first_counter1_1 = tlMasterXbar_monitor_1_a_first_counter_1 -10'h1; 
    wire tlMasterXbar_monitor_1_a_first_1 = tlMasterXbar_monitor_1_a_first_counter_1 ==10'h0; 
    wire[26:0] tlMasterXbar_monitor_1__d_first_beats1_decode_T_5 =27'hFFF<< tlMasterXbar_monitor_1__GEN_0 ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_beats1_decode_1 =~( tlMasterXbar_monitor_1__d_first_beats1_decode_T_5 [11:2]); 
    wire[9:0] tlMasterXbar_monitor_1_d_first_beats1_1 = tlMasterXbar_monitor_1_d_first_beats1_opdata_1  ?  tlMasterXbar_monitor_1_d_first_beats1_decode_1 :10'h0; reg[9:0] tlMasterXbar_monitor_1_d_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_counter1_1 = tlMasterXbar_monitor_1_d_first_counter_1 -10'h1; 
    wire tlMasterXbar_monitor_1_d_first_1 = tlMasterXbar_monitor_1_d_first_counter_1 ==10'h0; 
    wire tlMasterXbar_monitor_1_d_first_last_1 = tlMasterXbar_monitor_1_d_first_counter_1 ==10'h1| tlMasterXbar_monitor_1_d_first_beats1_1 ==10'h0; 
    wire tlMasterXbar_monitor_1_d_first_done_1 = tlMasterXbar_monitor_1_d_first_last_1 & tlMasterXbar_monitor_1_io_in_d_valid ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_count_1 = tlMasterXbar_monitor_1_d_first_beats1_1 &~ tlMasterXbar_monitor_1_d_first_counter1_1 ; 
    wire[3:0] tlMasterXbar_monitor_1_a_opcode_lookup ={1'h0, tlMasterXbar_monitor_1_inflight_opcodes [3:1]}; 
    wire[7:0] tlMasterXbar_monitor_1_a_size_lookup ={1'h0, tlMasterXbar_monitor_1_inflight_sizes [7:1]}; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_T_1 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_a_first_1 ; 
    wire tlMasterXbar_monitor_1_a_set_wo_ready ; 
  assign  tlMasterXbar_monitor_1_a_set_wo_ready = tlMasterXbar_monitor_1__same_cycle_resp_T_1 ; 
    wire tlMasterXbar_monitor_1_same_cycle_resp ; 
  assign  tlMasterXbar_monitor_1_same_cycle_resp = tlMasterXbar_monitor_1__same_cycle_resp_T_1 ; 
    wire tlMasterXbar_monitor_1_a_set = tlMasterXbar_monitor_1__a_first_T_1 & tlMasterXbar_monitor_1_a_first_1 ; 
    wire[3:0] tlMasterXbar_monitor_1_a_opcodes_set_interm = tlMasterXbar_monitor_1_a_set  ? 4'h9:4'h0; 
    wire[4:0] tlMasterXbar_monitor_1_a_sizes_set_interm = tlMasterXbar_monitor_1_a_set  ? 5'hD:5'h0; 
    wire[3:0] tlMasterXbar_monitor_1_a_opcodes_set = tlMasterXbar_monitor_1_a_set  ?  tlMasterXbar_monitor_1_a_opcodes_set_interm :4'h0; 
    wire[7:0] tlMasterXbar_monitor_1_a_sizes_set = tlMasterXbar_monitor_1_a_set  ? {3'h0, tlMasterXbar_monitor_1_a_sizes_set_interm }:8'h0; 
    wire tlMasterXbar_monitor_1__GEN_1 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_1 ; 
    wire tlMasterXbar_monitor_1__GEN_2 = tlMasterXbar_monitor_1__GEN_1 &~ tlMasterXbar_monitor_1_d_release_ack ; 
    wire tlMasterXbar_monitor_1_d_clr ; 
  assign  tlMasterXbar_monitor_1_d_clr = tlMasterXbar_monitor_1__GEN_2 ; 
    wire tlMasterXbar_monitor_1_d_clr_wo_ready ; 
  assign  tlMasterXbar_monitor_1_d_clr_wo_ready = tlMasterXbar_monitor_1__GEN_2 ; 
    wire[3:0] tlMasterXbar_monitor_1_d_opcodes_clr ={4{ tlMasterXbar_monitor_1__GEN_2 }}; 
    wire[7:0] tlMasterXbar_monitor_1_d_sizes_clr ={8{ tlMasterXbar_monitor_1__GEN_2 }}; reg[2:0] tlMasterXbar_monitor_1_casez_tmp ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_1_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h0;
              3 'b001: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h0;
              3 'b010: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h1;
              3 'b011: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h1;
              3 'b100: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h1;
              3 'b101: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h2;
              3 'b110: 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h4;
              default : 
                  tlMasterXbar_monitor_1_casez_tmp  =3'h4;endcase
         end
  reg[2:0] tlMasterXbar_monitor_1_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_1_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h0;
              3 'b001: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h0;
              3 'b010: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h1;
              3 'b011: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h1;
              3 'b100: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h1;
              3 'b101: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h2;
              3 'b110: 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h5;
              default : 
                  tlMasterXbar_monitor_1_casez_tmp_0  =3'h4;endcase
         end
  reg[31:0] tlMasterXbar_monitor_1_watchdog ; 
    reg tlMasterXbar_monitor_1_inflight_1 ; reg[3:0] tlMasterXbar_monitor_1_inflight_opcodes_1 ; reg[7:0] tlMasterXbar_monitor_1_inflight_sizes_1 ; 
    wire[26:0] tlMasterXbar_monitor_1__d_first_beats1_decode_T_9 =27'hFFF<< tlMasterXbar_monitor_1__GEN_0 ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_beats1_decode_2 =~( tlMasterXbar_monitor_1__d_first_beats1_decode_T_9 [11:2]); 
    wire[9:0] tlMasterXbar_monitor_1_d_first_beats1_2 = tlMasterXbar_monitor_1_d_first_beats1_opdata_2  ?  tlMasterXbar_monitor_1_d_first_beats1_decode_2 :10'h0; reg[9:0] tlMasterXbar_monitor_1_d_first_counter_2 ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_counter1_2 = tlMasterXbar_monitor_1_d_first_counter_2 -10'h1; 
    wire tlMasterXbar_monitor_1_d_first_2 = tlMasterXbar_monitor_1_d_first_counter_2 ==10'h0; 
    wire tlMasterXbar_monitor_1_d_first_last_2 = tlMasterXbar_monitor_1_d_first_counter_2 ==10'h1| tlMasterXbar_monitor_1_d_first_beats1_2 ==10'h0; 
    wire tlMasterXbar_monitor_1_d_first_done_2 = tlMasterXbar_monitor_1_d_first_last_2 & tlMasterXbar_monitor_1_io_in_d_valid ; 
    wire[9:0] tlMasterXbar_monitor_1_d_first_count_2 = tlMasterXbar_monitor_1_d_first_beats1_2 &~ tlMasterXbar_monitor_1_d_first_counter1_2 ; 
    wire[3:0] tlMasterXbar_monitor_1_c_opcode_lookup ={1'h0, tlMasterXbar_monitor_1_inflight_opcodes_1 [3:1]}; 
    wire[7:0] tlMasterXbar_monitor_1_c_size_lookup ={1'h0, tlMasterXbar_monitor_1_inflight_sizes_1 [7:1]}; 
    wire tlMasterXbar_monitor_1__GEN_3 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_2 & tlMasterXbar_monitor_1_d_release_ack_1 ; 
    wire tlMasterXbar_monitor_1_d_clr_1 ; 
  assign  tlMasterXbar_monitor_1_d_clr_1 = tlMasterXbar_monitor_1__GEN_3 ; 
    wire tlMasterXbar_monitor_1_d_clr_wo_ready_1 ; 
  assign  tlMasterXbar_monitor_1_d_clr_wo_ready_1 = tlMasterXbar_monitor_1__GEN_3 ; 
    wire[3:0] tlMasterXbar_monitor_1_d_opcodes_clr_1 ={4{ tlMasterXbar_monitor_1__GEN_3 }}; 
    wire[7:0] tlMasterXbar_monitor_1_d_sizes_clr_1 ={8{ tlMasterXbar_monitor_1__GEN_3 }}; reg[31:0] tlMasterXbar_monitor_1_watchdog_1 ; 
    wire tlMasterXbar_monitor_1__GEN_4 = tlMasterXbar_monitor_1_io_in_a_valid &~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_5 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1__GEN &~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_6 = tlMasterXbar_monitor_1_io_in_d_bits_size [3:1]==3'h0; 
    wire tlMasterXbar_monitor_1__GEN_7 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h4&~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_8 = tlMasterXbar_monitor_1_io_in_d_bits_param ==2'h2; 
    wire tlMasterXbar_monitor_1__GEN_9 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h5&~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_10 =~ tlMasterXbar_monitor_1_io_in_d_bits_denied | tlMasterXbar_monitor_1_io_in_d_bits_corrupt ; 
    wire tlMasterXbar_monitor_1__GEN_11 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h0&~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_12 = tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor_1__GEN_13 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1__GEN_12 &~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_14 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h2&~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_15 = tlMasterXbar_monitor_1_io_in_d_valid &~ tlMasterXbar_monitor_1_d_first &~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_16 = tlMasterXbar_monitor_1__GEN_2 & tlMasterXbar_monitor_1_same_cycle_resp &~ tlMasterXbar_monitor_1_reset ; 
    wire tlMasterXbar_monitor_1__GEN_17 = tlMasterXbar_monitor_1__GEN_2 &~ tlMasterXbar_monitor_1_same_cycle_resp &~ tlMasterXbar_monitor_1_reset ; 
    wire[7:0] tlMasterXbar_monitor_1__GEN_18 ={4'h0, tlMasterXbar_monitor_1_io_in_d_bits_size }; 
    wire tlMasterXbar_monitor_1__GEN_19 = tlMasterXbar_monitor_1__GEN_3 &~ tlMasterXbar_monitor_1_reset ; 
  always @( posedge  tlMasterXbar_monitor_1_clock )
         begin 
             if ( tlMasterXbar_monitor_1__GEN_4 &~({ tlMasterXbar_monitor_1_io_in_a_bits_address [31:14],~( tlMasterXbar_monitor_1_io_in_a_bits_address [13:12])}==20'h0| tlMasterXbar_monitor_1_io_in_a_bits_address [31:12]==20'h0|{ tlMasterXbar_monitor_1_io_in_a_bits_address [31:17],~( tlMasterXbar_monitor_1_io_in_a_bits_address [16])}==16'h0|{ tlMasterXbar_monitor_1_io_in_a_bits_address [31:26], tlMasterXbar_monitor_1_io_in_a_bits_address [25:16]^10'h200}==16'h0|{ tlMasterXbar_monitor_1_io_in_a_bits_address [31:28],~( tlMasterXbar_monitor_1_io_in_a_bits_address [27:26])}==6'h0|{ tlMasterXbar_monitor_1_io_in_a_bits_address [31],~( tlMasterXbar_monitor_1_io_in_a_bits_address [30:29])}==3'h0| tlMasterXbar_monitor_1_io_in_a_bits_address [31:14]==18'h20000))
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_4 &~ tlMasterXbar_monitor_1_is_aligned )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_io_in_d_valid &~ tlMasterXbar_monitor_1_reset &(& tlMasterXbar_monitor_1_io_in_d_bits_opcode ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_5 & tlMasterXbar_monitor_1__GEN_6 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_5 &(| tlMasterXbar_monitor_1_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_5 & tlMasterXbar_monitor_1_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_5 & tlMasterXbar_monitor_1_io_in_d_bits_denied )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_7 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_7 & tlMasterXbar_monitor_1__GEN_6 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_7 &(& tlMasterXbar_monitor_1_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_7 & tlMasterXbar_monitor_1__GEN_8 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_7 & tlMasterXbar_monitor_1_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_9 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_9 & tlMasterXbar_monitor_1__GEN_6 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_9 &(& tlMasterXbar_monitor_1_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_9 & tlMasterXbar_monitor_1__GEN_8 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_9 &~ tlMasterXbar_monitor_1__GEN_10 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_11 &(| tlMasterXbar_monitor_1_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_11 & tlMasterXbar_monitor_1_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_13 &(| tlMasterXbar_monitor_1_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_13 &~ tlMasterXbar_monitor_1__GEN_10 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_14 &(| tlMasterXbar_monitor_1_io_in_d_bits_param ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_14 & tlMasterXbar_monitor_1_io_in_d_bits_corrupt )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_io_in_a_valid &~ tlMasterXbar_monitor_1_a_first &~ tlMasterXbar_monitor_1_reset & tlMasterXbar_monitor_1_io_in_a_bits_address != tlMasterXbar_monitor_1_address )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_15 & tlMasterXbar_monitor_1_io_in_d_bits_opcode != tlMasterXbar_monitor_1_opcode_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_15 & tlMasterXbar_monitor_1_io_in_d_bits_param != tlMasterXbar_monitor_1_param_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_15 & tlMasterXbar_monitor_1_io_in_d_bits_size != tlMasterXbar_monitor_1_size_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_15 & tlMasterXbar_monitor_1_io_in_d_bits_sink != tlMasterXbar_monitor_1_sink )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_15 & tlMasterXbar_monitor_1_io_in_d_bits_denied != tlMasterXbar_monitor_1_denied )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_a_set &~ tlMasterXbar_monitor_1_reset & tlMasterXbar_monitor_1_inflight )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_2 &~ tlMasterXbar_monitor_1_reset &~( tlMasterXbar_monitor_1_inflight | tlMasterXbar_monitor_1_same_cycle_resp ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_16 &~ tlMasterXbar_monitor_1__GEN_12 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_16 & tlMasterXbar_monitor_1_io_in_d_bits_size !=4'h6)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_17 &~( tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_casez_tmp | tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_casez_tmp_0 ))
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_17 & tlMasterXbar_monitor_1__GEN_18 != tlMasterXbar_monitor_1_a_size_lookup )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_1 & tlMasterXbar_monitor_1_a_first_1 & tlMasterXbar_monitor_1_io_in_a_valid &~ tlMasterXbar_monitor_1_d_release_ack &~ tlMasterXbar_monitor_1_reset &~ tlMasterXbar_monitor_1_io_in_a_ready )
                 begin 
                     if (1)$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_monitor_1_reset &~( tlMasterXbar_monitor_1_a_set_wo_ready != tlMasterXbar_monitor_1_d_clr_wo_ready |~ tlMasterXbar_monitor_1_a_set_wo_ready ))
                 begin 
                     if (1)$error("Assertion failed: 'A' and 'D' concurrent, despite minlatency 4 (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_monitor_1_reset &~(~ tlMasterXbar_monitor_1_inflight | tlMasterXbar_monitor_1__plusarg_reader_out ==32'h0| tlMasterXbar_monitor_1_watchdog < tlMasterXbar_monitor_1__plusarg_reader_out ))
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_19 &~ tlMasterXbar_monitor_1_inflight_1 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_19 & tlMasterXbar_monitor_1__GEN_18 != tlMasterXbar_monitor_1_c_size_lookup )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (~ tlMasterXbar_monitor_1_reset &~(~ tlMasterXbar_monitor_1_inflight_1 | tlMasterXbar_monitor_1__plusarg_reader_1_out ==32'h0| tlMasterXbar_monitor_1_watchdog_1 < tlMasterXbar_monitor_1__plusarg_reader_1_out ))
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
         end
  always @( posedge  tlMasterXbar_monitor_1_clock )
         begin 
             if ( tlMasterXbar_monitor_1_reset )
                 begin  
                     tlMasterXbar_monitor_1_a_first_counter  <=10'h0; 
                     tlMasterXbar_monitor_1_d_first_counter  <=10'h0; 
                     tlMasterXbar_monitor_1_inflight  <=1'h0; 
                     tlMasterXbar_monitor_1_inflight_opcodes  <=4'h0; 
                     tlMasterXbar_monitor_1_inflight_sizes  <=8'h0; 
                     tlMasterXbar_monitor_1_a_first_counter_1  <=10'h0; 
                     tlMasterXbar_monitor_1_d_first_counter_1  <=10'h0; 
                     tlMasterXbar_monitor_1_watchdog  <=32'h0; 
                     tlMasterXbar_monitor_1_inflight_1  <=1'h0; 
                     tlMasterXbar_monitor_1_inflight_opcodes_1  <=4'h0; 
                     tlMasterXbar_monitor_1_inflight_sizes_1  <=8'h0; 
                     tlMasterXbar_monitor_1_d_first_counter_2  <=10'h0; 
                     tlMasterXbar_monitor_1_watchdog_1  <=32'h0;
                 end 
              else 
                 begin 
                     if ( tlMasterXbar_monitor_1__a_first_T_1 )
                         begin 
                             if ( tlMasterXbar_monitor_1_a_first ) 
                                 tlMasterXbar_monitor_1_a_first_counter  <=10'h0;
                              else  
                                 tlMasterXbar_monitor_1_a_first_counter  <= tlMasterXbar_monitor_1_a_first_counter1 ;
                             if ( tlMasterXbar_monitor_1_a_first_1 ) 
                                 tlMasterXbar_monitor_1_a_first_counter_1  <=10'h0;
                              else  
                                 tlMasterXbar_monitor_1_a_first_counter_1  <= tlMasterXbar_monitor_1_a_first_counter1_1 ;
                         end 
                     if ( tlMasterXbar_monitor_1_io_in_d_valid )
                         begin 
                             if ( tlMasterXbar_monitor_1_d_first ) 
                                 tlMasterXbar_monitor_1_d_first_counter  <= tlMasterXbar_monitor_1_d_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_1_d_first_counter  <= tlMasterXbar_monitor_1_d_first_counter1 ;
                             if ( tlMasterXbar_monitor_1_d_first_1 ) 
                                 tlMasterXbar_monitor_1_d_first_counter_1  <= tlMasterXbar_monitor_1_d_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_1_d_first_counter_1  <= tlMasterXbar_monitor_1_d_first_counter1_1 ;
                             if ( tlMasterXbar_monitor_1_d_first_2 ) 
                                 tlMasterXbar_monitor_1_d_first_counter_2  <= tlMasterXbar_monitor_1_d_first_beats1_2 ;
                              else  
                                 tlMasterXbar_monitor_1_d_first_counter_2  <= tlMasterXbar_monitor_1_d_first_counter1_2 ; 
                             tlMasterXbar_monitor_1_watchdog_1  <=32'h0;
                         end 
                      else  
                         tlMasterXbar_monitor_1_watchdog_1  <= tlMasterXbar_monitor_1_watchdog_1 +32'h1; 
                     tlMasterXbar_monitor_1_inflight  <=( tlMasterXbar_monitor_1_inflight | tlMasterXbar_monitor_1_a_set )&~ tlMasterXbar_monitor_1_d_clr ; 
                     tlMasterXbar_monitor_1_inflight_opcodes  <=( tlMasterXbar_monitor_1_inflight_opcodes | tlMasterXbar_monitor_1_a_opcodes_set )&~ tlMasterXbar_monitor_1_d_opcodes_clr ; 
                     tlMasterXbar_monitor_1_inflight_sizes  <=( tlMasterXbar_monitor_1_inflight_sizes | tlMasterXbar_monitor_1_a_sizes_set )&~ tlMasterXbar_monitor_1_d_sizes_clr ;
                     if ( tlMasterXbar_monitor_1__a_first_T_1 | tlMasterXbar_monitor_1_io_in_d_valid ) 
                         tlMasterXbar_monitor_1_watchdog  <=32'h0;
                      else  
                         tlMasterXbar_monitor_1_watchdog  <= tlMasterXbar_monitor_1_watchdog +32'h1; 
                     tlMasterXbar_monitor_1_inflight_1  <= tlMasterXbar_monitor_1_inflight_1 &~ tlMasterXbar_monitor_1_d_clr_1 ; 
                     tlMasterXbar_monitor_1_inflight_opcodes_1  <= tlMasterXbar_monitor_1_inflight_opcodes_1 &~ tlMasterXbar_monitor_1_d_opcodes_clr_1 ; 
                     tlMasterXbar_monitor_1_inflight_sizes_1  <= tlMasterXbar_monitor_1_inflight_sizes_1 &~ tlMasterXbar_monitor_1_d_sizes_clr_1 ;
                 end 
             if ( tlMasterXbar_monitor_1__a_first_T_1 & tlMasterXbar_monitor_1_a_first ) 
                 tlMasterXbar_monitor_1_address  <= tlMasterXbar_monitor_1_io_in_a_bits_address ;
             if ( tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first )
                 begin  
                     tlMasterXbar_monitor_1_opcode_1  <= tlMasterXbar_monitor_1_io_in_d_bits_opcode ; 
                     tlMasterXbar_monitor_1_param_1  <= tlMasterXbar_monitor_1_io_in_d_bits_param ; 
                     tlMasterXbar_monitor_1_size_1  <= tlMasterXbar_monitor_1_io_in_d_bits_size ; 
                     tlMasterXbar_monitor_1_sink  <= tlMasterXbar_monitor_1_io_in_d_bits_sink ; 
                     tlMasterXbar_monitor_1_denied  <= tlMasterXbar_monitor_1_io_in_d_bits_denied ;
                 end 
         end
    plusarg_reader  #(. tlMasterXbar_monitor_1_DEFAULT (0),. tlMasterXbar_monitor_1_FORMAT ("tilelink_timeout=%d"),. tlMasterXbar_monitor_1_WIDTH (32)) tlMasterXbar_monitor_1_plusarg_reader (. out ( tlMasterXbar_monitor_1__plusarg_reader_out ));  
    plusarg_reader  #(. tlMasterXbar_monitor_1_DEFAULT (0),. tlMasterXbar_monitor_1_FORMAT ("tilelink_timeout=%d"),. tlMasterXbar_monitor_1_WIDTH (32)) tlMasterXbar_monitor_1_plusarg_reader_1 (. out ( tlMasterXbar_monitor_1__plusarg_reader_1_out ));
    assign tlMasterXbar_monitor_1_clock = tlMasterXbar_clock;
    assign tlMasterXbar_monitor_1_reset = tlMasterXbar_reset;
    assign tlMasterXbar_monitor_1_io_in_a_ready = tlMasterXbar_nodeIn_1_a_ready;
    assign tlMasterXbar_monitor_1_io_in_a_valid = tlMasterXbar_nodeIn_1_a_valid;
    assign tlMasterXbar_monitor_1_io_in_a_bits_address = tlMasterXbar_nodeIn_1_a_bits_address;
    assign tlMasterXbar_monitor_1_io_in_d_valid = tlMasterXbar_nodeIn_1_d_valid;
    assign tlMasterXbar_monitor_1_io_in_d_bits_opcode = tlMasterXbar_nodeIn_1_d_bits_opcode;
    assign tlMasterXbar_monitor_1_io_in_d_bits_param = tlMasterXbar_nodeIn_1_d_bits_param;
    assign tlMasterXbar_monitor_1_io_in_d_bits_size = tlMasterXbar_nodeIn_1_d_bits_size;
    assign tlMasterXbar_monitor_1_io_in_d_bits_sink = tlMasterXbar_nodeIn_1_d_bits_sink;
    assign tlMasterXbar_monitor_1_io_in_d_bits_denied = tlMasterXbar_nodeIn_1_d_bits_denied;
    assign tlMasterXbar_monitor_1_io_in_d_bits_corrupt = tlMasterXbar_nodeIn_1_d_bits_corrupt;
     
  assign  tlMasterXbar_auto_in_1_a_ready = tlMasterXbar_nodeIn_1_a_ready ; 
  assign  tlMasterXbar_auto_in_1_d_valid = tlMasterXbar_nodeIn_1_d_valid ; 
  assign  tlMasterXbar_auto_in_1_d_bits_opcode = tlMasterXbar_nodeIn_1_d_bits_opcode ; 
  assign  tlMasterXbar_auto_in_1_d_bits_param = tlMasterXbar_nodeIn_1_d_bits_param ; 
  assign  tlMasterXbar_auto_in_1_d_bits_size = tlMasterXbar_nodeIn_1_d_bits_size ; 
  assign  tlMasterXbar_auto_in_1_d_bits_sink = tlMasterXbar_nodeIn_1_d_bits_sink ; 
  assign  tlMasterXbar_auto_in_1_d_bits_denied = tlMasterXbar_nodeIn_1_d_bits_denied ; 
  assign  tlMasterXbar_auto_in_1_d_bits_data = tlMasterXbar_nodeIn_1_d_bits_data ; 
  assign  tlMasterXbar_auto_in_1_d_bits_corrupt = tlMasterXbar_nodeIn_1_d_bits_corrupt ; 
  assign  tlMasterXbar_auto_in_0_a_ready = tlMasterXbar_nodeIn_a_ready ; 
  assign  tlMasterXbar_auto_in_0_d_valid = tlMasterXbar_nodeIn_d_valid ; 
  assign  tlMasterXbar_auto_in_0_d_bits_opcode = tlMasterXbar_nodeIn_d_bits_opcode ; 
  assign  tlMasterXbar_auto_in_0_d_bits_param = tlMasterXbar_nodeIn_d_bits_param ; 
  assign  tlMasterXbar_auto_in_0_d_bits_size = tlMasterXbar_nodeIn_d_bits_size ; 
  assign  tlMasterXbar_auto_in_0_d_bits_sink = tlMasterXbar_nodeIn_d_bits_sink ; 
  assign  tlMasterXbar_auto_in_0_d_bits_denied = tlMasterXbar_nodeIn_d_bits_denied ; 
  assign  tlMasterXbar_auto_in_0_d_bits_data = tlMasterXbar_nodeIn_d_bits_data ; 
  assign  tlMasterXbar_auto_in_0_d_bits_corrupt = tlMasterXbar_nodeIn_d_bits_corrupt ; 
  assign  tlMasterXbar_auto_out_a_valid = tlMasterXbar_nodeOut_a_valid ; 
  assign  tlMasterXbar_auto_out_a_bits_opcode = tlMasterXbar_nodeOut_a_bits_opcode ; 
  assign  tlMasterXbar_auto_out_a_bits_param = tlMasterXbar_nodeOut_a_bits_param ; 
  assign  tlMasterXbar_auto_out_a_bits_size = tlMasterXbar_nodeOut_a_bits_size ; 
  assign  tlMasterXbar_auto_out_a_bits_source = tlMasterXbar_nodeOut_a_bits_source ; 
  assign  tlMasterXbar_auto_out_a_bits_address = tlMasterXbar_nodeOut_a_bits_address ; 
  assign  tlMasterXbar_auto_out_a_bits_mask = tlMasterXbar_nodeOut_a_bits_mask ; 
  assign  tlMasterXbar_auto_out_a_bits_data = tlMasterXbar_nodeOut_a_bits_data ; 
  assign  tlMasterXbar_auto_out_d_ready = tlMasterXbar_nodeOut_d_ready ;
    assign tlMasterXbar_clock = clock;
    assign tlMasterXbar_reset = reset;
    assign widget_1_nodeOut_a_ready = tlMasterXbar_auto_in_1_a_ready;
    assign tlMasterXbar_auto_in_1_a_valid = widget_1_nodeOut_a_valid;
    assign tlMasterXbar_auto_in_1_a_bits_address = widget_1_nodeOut_a_bits_address;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_readalloc = widget_1_nodeOut_a_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_writealloc = widget_1_nodeOut_a_bits_user_amba_prot_writealloc;
    assign widget_1_nodeOut_d_valid = tlMasterXbar_auto_in_1_d_valid;
    assign widget_1_nodeOut_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode;
    assign widget_1_nodeOut_d_bits_param = tlMasterXbar_auto_in_1_d_bits_param;
    assign widget_1_nodeOut_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size;
    assign widget_1_nodeOut_d_bits_sink = tlMasterXbar_auto_in_1_d_bits_sink;
    assign widget_1_nodeOut_d_bits_denied = tlMasterXbar_auto_in_1_d_bits_denied;
    assign widget_1_nodeOut_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data;
    assign widget_1_nodeOut_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt;
    assign widget_nodeOut_a_ready = tlMasterXbar_auto_in_0_a_ready;
    assign tlMasterXbar_auto_in_0_a_valid = widget_nodeOut_a_valid;
    assign tlMasterXbar_auto_in_0_a_bits_opcode = widget_nodeOut_a_bits_opcode;
    assign tlMasterXbar_auto_in_0_a_bits_param = widget_nodeOut_a_bits_param;
    assign tlMasterXbar_auto_in_0_a_bits_size = widget_nodeOut_a_bits_size;
    assign tlMasterXbar_auto_in_0_a_bits_address = widget_nodeOut_a_bits_address;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_bufferable = widget_nodeOut_a_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_modifiable = widget_nodeOut_a_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_readalloc = widget_nodeOut_a_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_writealloc = widget_nodeOut_a_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_privileged = widget_nodeOut_a_bits_user_amba_prot_privileged;
    assign tlMasterXbar_auto_in_0_a_bits_mask = widget_nodeOut_a_bits_mask;
    assign tlMasterXbar_auto_in_0_a_bits_data = widget_nodeOut_a_bits_data;
    assign tlMasterXbar_auto_in_0_d_ready = widget_nodeOut_d_ready;
    assign widget_nodeOut_d_valid = tlMasterXbar_auto_in_0_d_valid;
    assign widget_nodeOut_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode;
    assign widget_nodeOut_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param;
    assign widget_nodeOut_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size;
    assign widget_nodeOut_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink;
    assign widget_nodeOut_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied;
    assign widget_nodeOut_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data;
    assign widget_nodeOut_d_bits_corrupt = tlMasterXbar_auto_in_0_d_bits_corrupt;
    assign tlMasterXbar_auto_out_a_ready = tlOtherMastersNodeIn_a_ready;
    assign tlOtherMastersNodeIn_a_valid = tlMasterXbar_auto_out_a_valid;
    assign tlOtherMastersNodeIn_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode;
    assign tlOtherMastersNodeIn_a_bits_param = tlMasterXbar_auto_out_a_bits_param;
    assign tlOtherMastersNodeIn_a_bits_size = tlMasterXbar_auto_out_a_bits_size;
    assign tlOtherMastersNodeIn_a_bits_source = tlMasterXbar_auto_out_a_bits_source;
    assign tlOtherMastersNodeIn_a_bits_address = tlMasterXbar_auto_out_a_bits_address;
    assign tlOtherMastersNodeIn_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask;
    assign tlOtherMastersNodeIn_a_bits_data = tlMasterXbar_auto_out_a_bits_data;
    assign tlOtherMastersNodeIn_d_ready = tlMasterXbar_auto_out_d_ready;
    assign tlMasterXbar_auto_out_d_valid = tlOtherMastersNodeIn_d_valid;
    assign tlMasterXbar_auto_out_d_bits_opcode = tlOtherMastersNodeIn_d_bits_opcode;
    assign tlMasterXbar_auto_out_d_bits_param = tlOtherMastersNodeIn_d_bits_param;
    assign tlMasterXbar_auto_out_d_bits_size = tlOtherMastersNodeIn_d_bits_size;
    assign tlMasterXbar_auto_out_d_bits_source = tlOtherMastersNodeIn_d_bits_source;
    assign tlMasterXbar_auto_out_d_bits_sink = tlOtherMastersNodeIn_d_bits_sink;
    assign tlMasterXbar_auto_out_d_bits_denied = tlOtherMastersNodeIn_d_bits_denied;
    assign tlMasterXbar_auto_out_d_bits_data = tlOtherMastersNodeIn_d_bits_data;
    assign tlMasterXbar_auto_out_d_bits_corrupt = tlOtherMastersNodeIn_d_bits_corrupt;
    
  wire intXbar_auto_int_in_2_0;
    wire intXbar_auto_int_in_1_0;
    wire intXbar_auto_int_in_1_1;
    wire intXbar_auto_int_in_0_0;
    wire intXbar_auto_int_out_0;
    wire intXbar_auto_int_out_1;
    wire intXbar_auto_int_out_2;
    wire intXbar_auto_int_out_3;

    wire intXbar_intnodeIn_0 = intXbar_auto_int_in_0_0 ; 
    wire intXbar_intnodeIn_1_0 = intXbar_auto_int_in_1_0 ; 
    wire intXbar_intnodeIn_1_1 = intXbar_auto_int_in_1_1 ; 
    wire intXbar_intnodeIn_2_0 = intXbar_auto_int_in_2_0 ; 
    wire intXbar_intnodeOut_0 = intXbar_intnodeIn_0 ; 
    wire intXbar_intnodeOut_1 = intXbar_intnodeIn_1_0 ; 
    wire intXbar_intnodeOut_2 = intXbar_intnodeIn_1_1 ; 
    wire intXbar_intnodeOut_3 = intXbar_intnodeIn_2_0 ; 
  assign  intXbar_auto_int_out_0 = intXbar_intnodeOut_0 ; 
  assign  intXbar_auto_int_out_1 = intXbar_intnodeOut_1 ; 
  assign  intXbar_auto_int_out_2 = intXbar_intnodeOut_2 ; 
  assign  intXbar_auto_int_out_3 = intXbar_intnodeOut_3 ;
    assign intXbar_auto_int_in_2_0 = x1_int_localOut_1_0;
    assign intXbar_auto_int_in_1_0 = x1_int_localOut_0;
    assign intXbar_auto_int_in_1_1 = x1_int_localOut_1;
    assign intXbar_auto_int_in_0_0 = int_localOut_0;
    assign intSinkNodeIn_0 = intXbar_auto_int_out_0;
    assign intSinkNodeIn_1 = intXbar_auto_int_out_1;
    assign intSinkNodeIn_2 = intXbar_auto_int_out_2;
    assign intSinkNodeIn_3 = intXbar_auto_int_out_3;
    
  wire dcache_clock;
    wire dcache_reset;
    wire dcache_auto_hart_id_sink_in;
    wire dcache_auto_out_a_ready;
    wire dcache_auto_out_a_valid;
    wire[2:0] dcache_auto_out_a_bits_opcode;
    wire[2:0] dcache_auto_out_a_bits_param;
    wire[3:0] dcache_auto_out_a_bits_size;
    wire[31:0] dcache_auto_out_a_bits_address;
    wire dcache_auto_out_a_bits_user_amba_prot_bufferable;
    wire dcache_auto_out_a_bits_user_amba_prot_modifiable;
    wire dcache_auto_out_a_bits_user_amba_prot_readalloc;
    wire dcache_auto_out_a_bits_user_amba_prot_writealloc;
    wire dcache_auto_out_a_bits_user_amba_prot_privileged;
    wire[3:0] dcache_auto_out_a_bits_mask;
    wire[31:0] dcache_auto_out_a_bits_data;
    wire dcache_auto_out_d_ready;
    wire dcache_auto_out_d_valid;
    wire[2:0] dcache_auto_out_d_bits_opcode;
    wire[1:0] dcache_auto_out_d_bits_param;
    wire[3:0] dcache_auto_out_d_bits_size;
    wire dcache_auto_out_d_bits_sink;
    wire dcache_auto_out_d_bits_denied;
    wire[31:0] dcache_auto_out_d_bits_data;
    wire dcache_auto_out_d_bits_corrupt;
    wire dcache_io_cpu_req_ready;
    wire dcache_io_cpu_req_valid;
    wire[31:0] dcache_io_cpu_req_bits_addr;
    wire[6:0] dcache_io_cpu_req_bits_tag;
    wire[4:0] dcache_io_cpu_req_bits_cmd;
    wire[1:0] dcache_io_cpu_req_bits_size;
    wire dcache_io_cpu_req_bits_signed;
    wire[1:0] dcache_io_cpu_req_bits_dprv;
    wire dcache_io_cpu_req_bits_dv;
    wire dcache_io_cpu_req_bits_phys;
    wire dcache_io_cpu_req_bits_no_xcpt;
    wire dcache_io_cpu_s1_kill;
    wire[31:0] dcache_io_cpu_s1_data_data;
    wire[3:0] dcache_io_cpu_s1_data_mask;
    wire dcache_io_cpu_s2_nack;
    wire dcache_io_cpu_resp_valid;
    wire[31:0] dcache_io_cpu_resp_bits_addr;
    wire[6:0] dcache_io_cpu_resp_bits_tag;
    wire[4:0] dcache_io_cpu_resp_bits_cmd;
    wire[1:0] dcache_io_cpu_resp_bits_size;
    wire dcache_io_cpu_resp_bits_signed;
    wire[1:0] dcache_io_cpu_resp_bits_dprv;
    wire dcache_io_cpu_resp_bits_dv;
    wire[31:0] dcache_io_cpu_resp_bits_data;
    wire[3:0] dcache_io_cpu_resp_bits_mask;
    wire dcache_io_cpu_resp_bits_replay;
    wire dcache_io_cpu_resp_bits_has_data;
    wire[31:0] dcache_io_cpu_resp_bits_data_word_bypass;
    wire[31:0] dcache_io_cpu_resp_bits_data_raw;
    wire[31:0] dcache_io_cpu_resp_bits_store_data;
    wire dcache_io_cpu_replay_next;
    wire dcache_io_cpu_s2_xcpt_ma_ld;
    wire dcache_io_cpu_s2_xcpt_ma_st;
    wire dcache_io_cpu_s2_xcpt_pf_ld;
    wire dcache_io_cpu_s2_xcpt_pf_st;
    wire dcache_io_cpu_s2_xcpt_ae_ld;
    wire dcache_io_cpu_s2_xcpt_ae_st;
    wire dcache_io_cpu_ordered;
    wire dcache_io_cpu_perf_grant;
    wire[19:0] dcache_io_ptw_req_bits_bits_addr;
    wire dcache_io_ptw_req_bits_bits_need_gpa;
    wire dcache_io_ptw_req_bits_bits_vstage1;
    wire dcache_io_ptw_req_bits_bits_stage2;
    wire dcache_io_ptw_resp_bits_ae_ptw;
    wire dcache_io_ptw_resp_bits_ae_final;
    wire dcache_io_ptw_resp_bits_pf;
    wire dcache_io_ptw_resp_bits_gf;
    wire dcache_io_ptw_resp_bits_hr;
    wire dcache_io_ptw_resp_bits_hw;
    wire dcache_io_ptw_resp_bits_hx;
    wire[43:0] dcache_io_ptw_resp_bits_pte_ppn;
    wire dcache_io_ptw_resp_bits_pte_d;
    wire dcache_io_ptw_resp_bits_pte_a;
    wire dcache_io_ptw_resp_bits_pte_g;
    wire dcache_io_ptw_resp_bits_pte_u;
    wire dcache_io_ptw_resp_bits_pte_x;
    wire dcache_io_ptw_resp_bits_pte_w;
    wire dcache_io_ptw_resp_bits_pte_r;
    wire dcache_io_ptw_resp_bits_pte_v;
    wire dcache_io_ptw_resp_bits_gpa_is_pte;
    wire dcache_io_ptw_status_debug;
    wire dcache_io_ptw_pmp_0_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_0_cfg_a;
    wire dcache_io_ptw_pmp_0_cfg_x;
    wire dcache_io_ptw_pmp_0_cfg_w;
    wire dcache_io_ptw_pmp_0_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_0_addr;
    wire[31:0] dcache_io_ptw_pmp_0_mask;
    wire dcache_io_ptw_pmp_1_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_1_cfg_a;
    wire dcache_io_ptw_pmp_1_cfg_x;
    wire dcache_io_ptw_pmp_1_cfg_w;
    wire dcache_io_ptw_pmp_1_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_1_addr;
    wire[31:0] dcache_io_ptw_pmp_1_mask;
    wire dcache_io_ptw_pmp_2_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_2_cfg_a;
    wire dcache_io_ptw_pmp_2_cfg_x;
    wire dcache_io_ptw_pmp_2_cfg_w;
    wire dcache_io_ptw_pmp_2_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_2_addr;
    wire[31:0] dcache_io_ptw_pmp_2_mask;
    wire dcache_io_ptw_pmp_3_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_3_cfg_a;
    wire dcache_io_ptw_pmp_3_cfg_x;
    wire dcache_io_ptw_pmp_3_cfg_w;
    wire dcache_io_ptw_pmp_3_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_3_addr;
    wire[31:0] dcache_io_ptw_pmp_3_mask;
    wire dcache_io_ptw_pmp_4_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_4_cfg_a;
    wire dcache_io_ptw_pmp_4_cfg_x;
    wire dcache_io_ptw_pmp_4_cfg_w;
    wire dcache_io_ptw_pmp_4_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_4_addr;
    wire[31:0] dcache_io_ptw_pmp_4_mask;
    wire dcache_io_ptw_pmp_5_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_5_cfg_a;
    wire dcache_io_ptw_pmp_5_cfg_x;
    wire dcache_io_ptw_pmp_5_cfg_w;
    wire dcache_io_ptw_pmp_5_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_5_addr;
    wire[31:0] dcache_io_ptw_pmp_5_mask;
    wire dcache_io_ptw_pmp_6_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_6_cfg_a;
    wire dcache_io_ptw_pmp_6_cfg_x;
    wire dcache_io_ptw_pmp_6_cfg_w;
    wire dcache_io_ptw_pmp_6_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_6_addr;
    wire[31:0] dcache_io_ptw_pmp_6_mask;
    wire dcache_io_ptw_pmp_7_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_7_cfg_a;
    wire dcache_io_ptw_pmp_7_cfg_x;
    wire dcache_io_ptw_pmp_7_cfg_w;
    wire dcache_io_ptw_pmp_7_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_7_addr;
    wire[31:0] dcache_io_ptw_pmp_7_mask;

    wire dcache__io_cpu_replay_next_output ; 
    wire dcache__io_cpu_s2_xcpt_ma_st_output ; 
    wire dcache__io_cpu_s2_xcpt_ma_ld_output ; 
    wire dcache__io_cpu_s2_xcpt_ae_st_output ; 
    wire dcache__io_cpu_s2_xcpt_ae_ld_output ; 
    wire dcache__io_cpu_s2_xcpt_pf_st_output ; 
    wire dcache__io_cpu_s2_xcpt_pf_ld_output ; 
    wire dcache__GEN ; 
    wire dcache_dataArb_io_in_1_valid ; 
    wire dcache_metaArb_io_in_3_valid ; 
    wire dcache_data_plaOutput ; 
    wire[3:0] dcache_dataArb_io_in_1_bits_eccMask ; 
    wire[13:0] dcache__dataArb_io_in_0_bits_wordMask_wordMask_T ; 
    wire dcache_dataArb_io_in_0_valid ; 
    wire dcache_metaArb_io_in_2_valid ; 
    wire[31:0] dcache_s1_all_data_ways_0 ; 
    wire[31:0] dcache_tl_d_data_encoded ; 
    wire[13:0] dcache_dataArb_io_in_3_bits_addr ; 
    wire[17:0] dcache__metaArb_io_in_5_bits_addr_T ; 
    wire dcache_dataArb_io_in_3_valid ; reg[1:0] dcache_s1_tlb_req_prv ; reg[4:0] dcache_s1_tlb_req_cmd ; reg[1:0] dcache_s1_tlb_req_size ; reg[31:0] dcache_s1_tlb_req_vaddr ; reg[1:0] dcache_s1_req_dprv ; reg[1:0] dcache_s1_req_size ; reg[4:0] dcache_s1_req_cmd ; reg[31:0] dcache_s1_req_addr ; 
    wire dcache_s0_req_phys ; 
    wire[31:0] dcache_s0_req_addr ; 
    wire[31:0] dcache_tl_out_a_bits_data ; 
    wire[3:0] dcache_tl_out_a_bits_mask ; 
    wire dcache_tl_out_a_bits_user_amba_prot_privileged ; 
    wire dcache_tl_out_a_bits_user_amba_prot_writealloc ; 
    wire dcache_tl_out_a_bits_user_amba_prot_readalloc ; 
    wire dcache_tl_out_a_bits_user_amba_prot_modifiable ; 
    wire dcache_tl_out_a_bits_user_amba_prot_bufferable ; 
    wire[31:0] dcache_tl_out_a_bits_address ; 
    wire[3:0] dcache_tl_out_a_bits_size ; 
    wire[2:0] dcache_tl_out_a_bits_param ; 
    wire[2:0] dcache_tl_out_a_bits_opcode ; 
    wire dcache_tl_out_a_valid ; 
    wire[31:0] dcache__amoalus_0_io_out_unmasked ; 
    wire dcache__lfsr_prng_io_out_0 ; 
    wire dcache__lfsr_prng_io_out_1 ; 
    wire dcache__lfsr_prng_io_out_2 ; 
    wire dcache__lfsr_prng_io_out_3 ; 
    wire dcache__lfsr_prng_io_out_4 ; 
    wire dcache__lfsr_prng_io_out_5 ; 
    wire dcache__lfsr_prng_io_out_6 ; 
    wire dcache__lfsr_prng_io_out_7 ; 
    wire dcache__lfsr_prng_io_out_8 ; 
    wire dcache__lfsr_prng_io_out_9 ; 
    wire dcache__lfsr_prng_io_out_10 ; 
    wire dcache__lfsr_prng_io_out_11 ; 
    wire dcache__lfsr_prng_io_out_12 ; 
    wire dcache__lfsr_prng_io_out_13 ; 
    wire dcache__lfsr_prng_io_out_14 ; 
    wire dcache__lfsr_prng_io_out_15 ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_c ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_c ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_c ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_c ; 
    wire dcache__pma_checker_entries_barrier_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_io_y_c ; 
    wire dcache__pma_checker_pmp_io_r ; 
    wire dcache__pma_checker_pmp_io_w ; 
    wire dcache__pma_checker_pmp_io_x ; 
    wire dcache__tlb_entries_barrier_5_io_y_u ; 
    wire dcache__tlb_entries_barrier_5_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_5_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_5_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_5_io_y_pf ; 
    wire dcache__tlb_entries_barrier_5_io_y_gf ; 
    wire dcache__tlb_entries_barrier_5_io_y_sw ; 
    wire dcache__tlb_entries_barrier_5_io_y_sx ; 
    wire dcache__tlb_entries_barrier_5_io_y_sr ; 
    wire dcache__tlb_entries_barrier_5_io_y_hw ; 
    wire dcache__tlb_entries_barrier_5_io_y_hx ; 
    wire dcache__tlb_entries_barrier_5_io_y_hr ; 
    wire dcache__tlb_entries_barrier_4_io_y_u ; 
    wire dcache__tlb_entries_barrier_4_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_4_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_4_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_4_io_y_pf ; 
    wire dcache__tlb_entries_barrier_4_io_y_gf ; 
    wire dcache__tlb_entries_barrier_4_io_y_sw ; 
    wire dcache__tlb_entries_barrier_4_io_y_sx ; 
    wire dcache__tlb_entries_barrier_4_io_y_sr ; 
    wire dcache__tlb_entries_barrier_4_io_y_hw ; 
    wire dcache__tlb_entries_barrier_4_io_y_hx ; 
    wire dcache__tlb_entries_barrier_4_io_y_hr ; 
    wire dcache__tlb_entries_barrier_4_io_y_pw ; 
    wire dcache__tlb_entries_barrier_4_io_y_px ; 
    wire dcache__tlb_entries_barrier_4_io_y_pr ; 
    wire dcache__tlb_entries_barrier_4_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_4_io_y_pal ; 
    wire dcache__tlb_entries_barrier_4_io_y_paa ; 
    wire dcache__tlb_entries_barrier_4_io_y_eff ; 
    wire dcache__tlb_entries_barrier_4_io_y_c ; 
    wire dcache__tlb_entries_barrier_3_io_y_u ; 
    wire dcache__tlb_entries_barrier_3_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_3_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_3_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_3_io_y_pf ; 
    wire dcache__tlb_entries_barrier_3_io_y_gf ; 
    wire dcache__tlb_entries_barrier_3_io_y_sw ; 
    wire dcache__tlb_entries_barrier_3_io_y_sx ; 
    wire dcache__tlb_entries_barrier_3_io_y_sr ; 
    wire dcache__tlb_entries_barrier_3_io_y_hw ; 
    wire dcache__tlb_entries_barrier_3_io_y_hx ; 
    wire dcache__tlb_entries_barrier_3_io_y_hr ; 
    wire dcache__tlb_entries_barrier_3_io_y_pw ; 
    wire dcache__tlb_entries_barrier_3_io_y_px ; 
    wire dcache__tlb_entries_barrier_3_io_y_pr ; 
    wire dcache__tlb_entries_barrier_3_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_3_io_y_pal ; 
    wire dcache__tlb_entries_barrier_3_io_y_paa ; 
    wire dcache__tlb_entries_barrier_3_io_y_eff ; 
    wire dcache__tlb_entries_barrier_3_io_y_c ; 
    wire dcache__tlb_entries_barrier_2_io_y_u ; 
    wire dcache__tlb_entries_barrier_2_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_2_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_2_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_2_io_y_pf ; 
    wire dcache__tlb_entries_barrier_2_io_y_gf ; 
    wire dcache__tlb_entries_barrier_2_io_y_sw ; 
    wire dcache__tlb_entries_barrier_2_io_y_sx ; 
    wire dcache__tlb_entries_barrier_2_io_y_sr ; 
    wire dcache__tlb_entries_barrier_2_io_y_hw ; 
    wire dcache__tlb_entries_barrier_2_io_y_hx ; 
    wire dcache__tlb_entries_barrier_2_io_y_hr ; 
    wire dcache__tlb_entries_barrier_2_io_y_pw ; 
    wire dcache__tlb_entries_barrier_2_io_y_px ; 
    wire dcache__tlb_entries_barrier_2_io_y_pr ; 
    wire dcache__tlb_entries_barrier_2_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_2_io_y_pal ; 
    wire dcache__tlb_entries_barrier_2_io_y_paa ; 
    wire dcache__tlb_entries_barrier_2_io_y_eff ; 
    wire dcache__tlb_entries_barrier_2_io_y_c ; 
    wire dcache__tlb_entries_barrier_1_io_y_u ; 
    wire dcache__tlb_entries_barrier_1_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_1_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_1_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_1_io_y_pf ; 
    wire dcache__tlb_entries_barrier_1_io_y_gf ; 
    wire dcache__tlb_entries_barrier_1_io_y_sw ; 
    wire dcache__tlb_entries_barrier_1_io_y_sx ; 
    wire dcache__tlb_entries_barrier_1_io_y_sr ; 
    wire dcache__tlb_entries_barrier_1_io_y_hw ; 
    wire dcache__tlb_entries_barrier_1_io_y_hx ; 
    wire dcache__tlb_entries_barrier_1_io_y_hr ; 
    wire dcache__tlb_entries_barrier_1_io_y_pw ; 
    wire dcache__tlb_entries_barrier_1_io_y_px ; 
    wire dcache__tlb_entries_barrier_1_io_y_pr ; 
    wire dcache__tlb_entries_barrier_1_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_1_io_y_pal ; 
    wire dcache__tlb_entries_barrier_1_io_y_paa ; 
    wire dcache__tlb_entries_barrier_1_io_y_eff ; 
    wire dcache__tlb_entries_barrier_1_io_y_c ; 
    wire dcache__tlb_entries_barrier_io_y_u ; 
    wire dcache__tlb_entries_barrier_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_io_y_pf ; 
    wire dcache__tlb_entries_barrier_io_y_gf ; 
    wire dcache__tlb_entries_barrier_io_y_sw ; 
    wire dcache__tlb_entries_barrier_io_y_sx ; 
    wire dcache__tlb_entries_barrier_io_y_sr ; 
    wire dcache__tlb_entries_barrier_io_y_hw ; 
    wire dcache__tlb_entries_barrier_io_y_hx ; 
    wire dcache__tlb_entries_barrier_io_y_hr ; 
    wire dcache__tlb_entries_barrier_io_y_pw ; 
    wire dcache__tlb_entries_barrier_io_y_px ; 
    wire dcache__tlb_entries_barrier_io_y_pr ; 
    wire dcache__tlb_entries_barrier_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_io_y_pal ; 
    wire dcache__tlb_entries_barrier_io_y_paa ; 
    wire dcache__tlb_entries_barrier_io_y_eff ; 
    wire dcache__tlb_entries_barrier_io_y_c ; 
    wire dcache__tlb_pmp_io_r ; 
    wire dcache__tlb_pmp_io_w ; 
    wire dcache__tlb_pmp_io_x ; 
    wire dcache_nodeOut_a_ready = dcache_auto_out_a_ready ; 
    wire dcache_nodeOut_d_valid = dcache_auto_out_d_valid ; 
    wire[2:0] dcache_nodeOut_d_bits_opcode = dcache_auto_out_d_bits_opcode ; 
    wire[1:0] dcache_nodeOut_d_bits_param = dcache_auto_out_d_bits_param ; 
    wire[3:0] dcache_nodeOut_d_bits_size = dcache_auto_out_d_bits_size ; 
    wire dcache_nodeOut_d_bits_sink = dcache_auto_out_d_bits_sink ; 
    wire dcache_nodeOut_d_bits_denied = dcache_auto_out_d_bits_denied ; 
    wire[31:0] dcache_nodeOut_d_bits_data = dcache_auto_out_d_bits_data ; 
    wire dcache_nodeOut_d_bits_corrupt = dcache_auto_out_d_bits_corrupt ; 
    wire dcache_hartIdSinkNodeOptIn = dcache_auto_hart_id_sink_in ; 
    wire dcache_tlb_newEntry_u = dcache_io_ptw_resp_bits_pte_u ; 
    wire dcache_tlb_newEntry_ae_ptw = dcache_io_ptw_resp_bits_ae_ptw ; 
    wire dcache_tlb_newEntry_ae_final = dcache_io_ptw_resp_bits_ae_final ; 
    wire dcache_tlb_newEntry_pf = dcache_io_ptw_resp_bits_pf ; 
    wire dcache_tlb_newEntry_gf = dcache_io_ptw_resp_bits_gf ; 
    wire dcache_tlb_newEntry_hw = dcache_io_ptw_resp_bits_hw ; 
    wire dcache_tlb_newEntry_hx = dcache_io_ptw_resp_bits_hx ; 
    wire dcache_tlb_newEntry_hr = dcache_io_ptw_resp_bits_hr ; 
    wire[6:0] dcache_s0_req_tag = dcache_io_cpu_req_bits_tag ; 
    wire[4:0] dcache_s0_req_cmd = dcache_io_cpu_req_bits_cmd ; 
    wire[1:0] dcache_s0_req_size = dcache_io_cpu_req_bits_size ; 
    wire dcache_s0_req_signed = dcache_io_cpu_req_bits_signed ; 
    wire[1:0] dcache_s0_req_dprv = dcache_io_cpu_req_bits_dprv ; 
    wire dcache_s0_req_dv = dcache_io_cpu_req_bits_dv ; 
    wire dcache_s0_req_no_xcpt = dcache_io_cpu_req_bits_no_xcpt ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_secure =1'h1; 
    wire dcache_metaArb_grant_1 =1'h1; 
    wire dcache_metaArb_grant_2 =1'h1; 
    wire dcache_tl_out_a_bits_user_amba_prot_secure =1'h1; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_secure =1'h1; 
    wire dcache_tl_out_c_bits_user_amba_prot_bufferable =1'h1; 
    wire dcache_tl_out_c_bits_user_amba_prot_modifiable =1'h1; 
    wire dcache_tl_out_c_bits_user_amba_prot_readalloc =1'h1; 
    wire dcache_tl_out_c_bits_user_amba_prot_writealloc =1'h1; 
    wire dcache_tl_out_c_bits_user_amba_prot_privileged =1'h1; 
    wire dcache_tl_out_c_bits_user_amba_prot_secure =1'h1; 
    wire dcache_a_sel =1'h1; 
    wire dcache_canAcceptCachedGrant =1'h1; 
    wire dcache_uncachedRespIdxOH =1'h1; 
    wire dcache_c_first =1'h1; 
    wire dcache_c_last =1'h1; 
    wire dcache_io_cpu_perf_release_first =1'h1; 
    wire dcache_io_cpu_perf_release_last =1'h1; 
    wire[24:0] dcache_pma_checker_special_entry_data_0_hi_hi =25'h0; 
    wire[24:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi =25'h0; 
    wire[24:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi =25'h0; 
    wire[24:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi =25'h0; 
    wire[24:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi =25'h0; 
    wire[24:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi =25'h0; 
    wire[1:0] dcache_hitState_meta_state =2'h3; 
    wire[5:0] dcache_tlb_real_hits =6'h0; 
    wire[5:0] dcache_tlb_stage1_bypass =6'h0; 
    wire[5:0] dcache_pma_checker_real_hits =6'h0; 
    wire[5:0] dcache_pma_checker_special_entry_data_0_hi_lo =6'h0; 
    wire[5:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo =6'h0; 
    wire[5:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo =6'h0; 
    wire[5:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo =6'h0; 
    wire[5:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo =6'h0; 
    wire[5:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo =6'h0; 
    wire[5:0] dcache_pma_checker_stage1_bypass =6'h0; 
    wire dcache_nodeOut_a_bits_source =1'h0; 
    wire dcache_nodeOut_a_bits_user_amba_prot_fetch =1'h0; 
    wire dcache_nodeOut_a_bits_corrupt =1'h0; 
    wire dcache_nodeOut_d_bits_source =1'h0; 
    wire dcache_mmioAddressPrefixSinkNodeOptIn =1'h0; 
    wire dcache_tlb_priv_v =1'h0; 
    wire dcache_tlb_satp_mode =1'h0; 
    wire dcache_tlb_stage1_en =1'h0; 
    wire dcache_tlb_vstage1_en =1'h0; 
    wire dcache_tlb_stage2_en =1'h0; 
    wire dcache_tlb_vm_enabled =1'h0; 
    wire dcache_tlb_vsatp_mode_mismatch =1'h0; 
    wire dcache_tlb_do_refill =1'h0; 
    wire dcache_tlb_cacheable =1'h0; 
    wire dcache_tlb_sector_hits_0 =1'h0; 
    wire dcache_tlb_superpage_hits_0 =1'h0; 
    wire dcache_tlb_superpage_hits_1 =1'h0; 
    wire dcache_tlb_superpage_hits_2 =1'h0; 
    wire dcache_tlb_superpage_hits_3 =1'h0; 
    wire dcache_tlb_hitsVec_0 =1'h0; 
    wire dcache_tlb_hitsVec_1 =1'h0; 
    wire dcache_tlb_hitsVec_2 =1'h0; 
    wire dcache_tlb_hitsVec_3 =1'h0; 
    wire dcache_tlb_hitsVec_4 =1'h0; 
    wire dcache_tlb_hitsVec_5 =1'h0; 
    wire dcache_tlb_refill_v =1'h0; 
    wire dcache_tlb_newEntry_ae_stage2 =1'h0; 
    wire dcache_tlb_newEntry_c =1'h0; 
    wire dcache_tlb_newEntry_fragmented_superpage =1'h0; 
    wire dcache_tlb_sum =1'h0; 
    wire dcache_tlb_mxr =1'h0; 
    wire dcache_tlb_cmd_readx =1'h0; 
    wire dcache_tlb_tlb_hit_if_not_gpa_miss =1'h0; 
    wire dcache_tlb_tlb_hit =1'h0; 
    wire dcache_tlb_tlb_miss =1'h0; 
    wire dcache_tlb_state_reg_left_subtree_state =1'h0; 
    wire dcache_tlb_state_reg_right_subtree_state =1'h0; 
    wire dcache_tlb_multipleHits_leftOne =1'h0; 
    wire dcache_tlb_multipleHits_leftOne_1 =1'h0; 
    wire dcache_tlb_multipleHits_rightOne =1'h0; 
    wire dcache_tlb_multipleHits_rightOne_1 =1'h0; 
    wire dcache_tlb_multipleHits_rightTwo =1'h0; 
    wire dcache_tlb_multipleHits_leftOne_2 =1'h0; 
    wire dcache_tlb_multipleHits_leftTwo =1'h0; 
    wire dcache_tlb_multipleHits_leftOne_3 =1'h0; 
    wire dcache_tlb_multipleHits_leftOne_4 =1'h0; 
    wire dcache_tlb_multipleHits_rightOne_2 =1'h0; 
    wire dcache_tlb_multipleHits_rightOne_3 =1'h0; 
    wire dcache_tlb_multipleHits_rightTwo_1 =1'h0; 
    wire dcache_tlb_multipleHits_rightOne_4 =1'h0; 
    wire dcache_tlb_multipleHits_rightTwo_2 =1'h0; 
    wire dcache_tlb_multipleHits =1'h0; 
    wire dcache_pma_checker_priv_v =1'h0; 
    wire dcache_pma_checker_satp_mode =1'h0; 
    wire dcache_pma_checker_stage1_en =1'h0; 
    wire dcache_pma_checker_vstage1_en =1'h0; 
    wire dcache_pma_checker_stage2_en =1'h0; 
    wire dcache_pma_checker_vm_enabled =1'h0; 
    wire dcache_pma_checker_vsatp_mode_mismatch =1'h0; 
    wire dcache_pma_checker_do_refill =1'h0; 
    wire dcache_pma_checker_invalidate_refill =1'h0; 
    wire dcache_pma_checker_cacheable =1'h0; 
    wire dcache_pma_checker_sector_hits_0 =1'h0; 
    wire dcache_pma_checker_superpage_hits_0 =1'h0; 
    wire dcache_pma_checker_superpage_hits_1 =1'h0; 
    wire dcache_pma_checker_superpage_hits_2 =1'h0; 
    wire dcache_pma_checker_superpage_hits_3 =1'h0; 
    wire dcache_pma_checker_hitsVec_0 =1'h0; 
    wire dcache_pma_checker_hitsVec_1 =1'h0; 
    wire dcache_pma_checker_hitsVec_2 =1'h0; 
    wire dcache_pma_checker_hitsVec_3 =1'h0; 
    wire dcache_pma_checker_hitsVec_4 =1'h0; 
    wire dcache_pma_checker_hitsVec_5 =1'h0; 
    wire dcache_pma_checker_refill_v =1'h0; 
    wire dcache_pma_checker_newEntry_u =1'h0; 
    wire dcache_pma_checker_newEntry_g =1'h0; 
    wire dcache_pma_checker_newEntry_ae_ptw =1'h0; 
    wire dcache_pma_checker_newEntry_ae_final =1'h0; 
    wire dcache_pma_checker_newEntry_ae_stage2 =1'h0; 
    wire dcache_pma_checker_newEntry_pf =1'h0; 
    wire dcache_pma_checker_newEntry_gf =1'h0; 
    wire dcache_pma_checker_newEntry_sw =1'h0; 
    wire dcache_pma_checker_newEntry_sx =1'h0; 
    wire dcache_pma_checker_newEntry_sr =1'h0; 
    wire dcache_pma_checker_newEntry_hw =1'h0; 
    wire dcache_pma_checker_newEntry_hx =1'h0; 
    wire dcache_pma_checker_newEntry_hr =1'h0; 
    wire dcache_pma_checker_newEntry_c =1'h0; 
    wire dcache_pma_checker_newEntry_fragmented_superpage =1'h0; 
    wire dcache_pma_checker_sum =1'h0; 
    wire dcache_pma_checker_mxr =1'h0; 
    wire dcache_pma_checker_cmd_readx =1'h0; 
    wire dcache_pma_checker_tlb_hit_if_not_gpa_miss =1'h0; 
    wire dcache_pma_checker_tlb_hit =1'h0; 
    wire dcache_pma_checker_tlb_miss =1'h0; 
    wire dcache_pma_checker_state_reg_left_subtree_state =1'h0; 
    wire dcache_pma_checker_state_reg_right_subtree_state =1'h0; 
    wire dcache_pma_checker_multipleHits_leftOne =1'h0; 
    wire dcache_pma_checker_multipleHits_leftOne_1 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightOne =1'h0; 
    wire dcache_pma_checker_multipleHits_rightOne_1 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightTwo =1'h0; 
    wire dcache_pma_checker_multipleHits_leftOne_2 =1'h0; 
    wire dcache_pma_checker_multipleHits_leftTwo =1'h0; 
    wire dcache_pma_checker_multipleHits_leftOne_3 =1'h0; 
    wire dcache_pma_checker_multipleHits_leftOne_4 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightOne_2 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightOne_3 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightTwo_1 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightOne_4 =1'h0; 
    wire dcache_pma_checker_multipleHits_rightTwo_2 =1'h0; 
    wire dcache_pma_checker_multipleHits =1'h0; 
    wire dcache_tl_out_a_bits_source =1'h0; 
    wire dcache_tl_out_a_bits_user_amba_prot_fetch =1'h0; 
    wire dcache_tl_out_a_bits_corrupt =1'h0; 
    wire dcache_nodeOut_a_deq_bits_source =1'h0; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_fetch =1'h0; 
    wire dcache_nodeOut_a_deq_bits_corrupt =1'h0; 
    wire dcache_tl_out_c_ready =1'h0; 
    wire dcache_tl_out_c_bits_user_amba_prot_fetch =1'h0; 
    wire dcache_tl_out_c_bits_corrupt =1'h0; 
    wire dcache_s0_req_no_alloc =1'h0; 
    wire dcache_s1_waw_hazard =1'h0; 
    wire dcache_inWriteback =1'h0; 
    wire dcache_s1_victim_way =1'h0; 
    wire dcache_releaseInFlight =1'h0; 
    wire dcache_s2_meta_error_uncorrectable =1'h0; 
    wire dcache_s2_meta_error =1'h0; 
    wire dcache_s2_store_merge =1'h0; 
    wire dcache_s2_data_error =1'h0; 
    wire dcache_s2_data_error_uncorrectable =1'h0; 
    wire dcache_s2_valid_data_error =1'h0; 
    wire dcache_s2_want_victimize =1'h0; 
    wire dcache_s2_cannot_victimize =1'h0; 
    wire dcache_s2_victimize =1'h0; 
    wire dcache_s2_lr =1'h0; 
    wire dcache_s2_sc =1'h0; 
    wire dcache_s2_sc_fail =1'h0; 
    wire dcache_s2_correct =1'h0; 
    wire dcache_s2_valid_correct =1'h0; 
    wire dcache_pstore1_merge_likely =1'h0; 
    wire dcache_pstore1_merge =1'h0; 
    wire dcache_pstore_drain_s2_kill =1'h0; 
    wire dcache_dataArb_io_in_0_valid_s2_kill =1'h0; 
    wire dcache_get_source =1'h0; 
    wire dcache_get_user_amba_prot_bufferable =1'h0; 
    wire dcache_get_user_amba_prot_modifiable =1'h0; 
    wire dcache_get_user_amba_prot_readalloc =1'h0; 
    wire dcache_get_user_amba_prot_writealloc =1'h0; 
    wire dcache_get_user_amba_prot_privileged =1'h0; 
    wire dcache_get_user_amba_prot_secure =1'h0; 
    wire dcache_get_user_amba_prot_fetch =1'h0; 
    wire dcache_get_corrupt =1'h0; 
    wire dcache_put_source =1'h0; 
    wire dcache_put_user_amba_prot_bufferable =1'h0; 
    wire dcache_put_user_amba_prot_modifiable =1'h0; 
    wire dcache_put_user_amba_prot_readalloc =1'h0; 
    wire dcache_put_user_amba_prot_writealloc =1'h0; 
    wire dcache_put_user_amba_prot_privileged =1'h0; 
    wire dcache_put_user_amba_prot_secure =1'h0; 
    wire dcache_put_user_amba_prot_fetch =1'h0; 
    wire dcache_put_corrupt =1'h0; 
    wire dcache_putpartial_source =1'h0; 
    wire dcache_putpartial_user_amba_prot_bufferable =1'h0; 
    wire dcache_putpartial_user_amba_prot_modifiable =1'h0; 
    wire dcache_putpartial_user_amba_prot_readalloc =1'h0; 
    wire dcache_putpartial_user_amba_prot_writealloc =1'h0; 
    wire dcache_putpartial_user_amba_prot_privileged =1'h0; 
    wire dcache_putpartial_user_amba_prot_secure =1'h0; 
    wire dcache_putpartial_user_amba_prot_fetch =1'h0; 
    wire dcache_putpartial_corrupt =1'h0; 
    wire dcache_atomics_a_source =1'h0; 
    wire dcache_atomics_a_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_corrupt =1'h0; 
    wire dcache_atomics_a_1_source =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_1_corrupt =1'h0; 
    wire dcache_atomics_a_2_source =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_2_corrupt =1'h0; 
    wire dcache_atomics_a_3_source =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_3_corrupt =1'h0; 
    wire dcache_atomics_a_4_source =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_4_corrupt =1'h0; 
    wire dcache_atomics_a_5_source =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_5_corrupt =1'h0; 
    wire dcache_atomics_a_6_source =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_6_corrupt =1'h0; 
    wire dcache_atomics_a_7_source =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_7_corrupt =1'h0; 
    wire dcache_atomics_a_8_source =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_8_corrupt =1'h0; 
    wire dcache_atomics_source =1'h0; 
    wire dcache_atomics_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_corrupt =1'h0; 
    wire dcache_grantIsCached =1'h0; 
    wire dcache_grantIsVoluntary =1'h0; 
    wire dcache_grantIsRefill =1'h0; 
    wire dcache_block_probe_for_pending_release_ack =1'h0; 
    wire dcache_beats1_opdata_1 =1'h0; 
    wire dcache_releaseDone =1'h0; 
    wire dcache_nackResponseMessage_source =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_bufferable =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_modifiable =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_readalloc =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_writealloc =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_privileged =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_secure =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_fetch =1'h0; 
    wire dcache_nackResponseMessage_corrupt =1'h0; 
    wire dcache_cleanReleaseMessage_source =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_bufferable =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_modifiable =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_readalloc =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_writealloc =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_privileged =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_secure =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_fetch =1'h0; 
    wire dcache_cleanReleaseMessage_corrupt =1'h0; 
    wire dcache_dirtyReleaseMessage_source =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_bufferable =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_modifiable =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_readalloc =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_writealloc =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_privileged =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_secure =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_fetch =1'h0; 
    wire dcache_dirtyReleaseMessage_corrupt =1'h0; 
    wire dcache_io_cpu_resp_bits_data_doZero =1'h0; 
    wire dcache_io_cpu_resp_bits_data_doZero_1 =1'h0; 
    wire dcache_flushDone =1'h0; 
    wire dcache_io_cpu_perf_release_beats1_opdata =1'h0; 
    wire dcache_io_cpu_perf_release_done =1'h0; 
    wire[9:0] dcache_counter1_1 =10'h3FF; 
    wire[9:0] dcache_io_cpu_perf_release_counter1 =10'h3FF; 
    wire[1:0] dcache_tlb_real_hits_lo_hi =2'h0; 
    wire[1:0] dcache_tlb_real_hits_hi_hi =2'h0; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_tlb_waddr =2'h0; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_tlb_idx =2'h0; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_real_hits_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_real_hits_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_hi_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_hi_lo_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_hi_lo_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_hi_hi_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_waddr =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_idx =2'h0; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo_lo =2'h0; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_lo_hi =2'h0; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_hi_hi =2'h0; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_lo_hi =2'h0; 
    wire[1:0] dcache_hitState_meta_1_state =2'h0; 
    wire[1:0] dcache_dummyMeta_meta_state =2'h0; 
    wire[1:0] dcache_dummyMeta_coh_state =2'h0; 
    wire[1:0] dcache_s2_valid_no_xcpt_lo_hi =2'h0; 
    wire[1:0] dcache_s2_meta_corrected_0_coh_state =2'h0; 
    wire[1:0] dcache_voluntaryNewCoh_state =2'h0; 
    wire[1:0] dcache_metaArb_io_in_1_bits_data_new_meta_coh_state =2'h0; 
    wire[1:0] dcache_metaArb_io_in_1_bits_data_new_meta_coh_meta_state =2'h0; 
    wire[1:0] dcache_metaArb_io_in_0_bits_data_meta_state =2'h0; 
    wire[1:0] dcache_metaArb_io_in_0_bits_data_meta_1_coh_state =2'h0; 
    wire[8:0] dcache_tlb_satp_asid =9'h0; 
    wire[8:0] dcache_pma_checker_satp_asid =9'h0; 
    wire[2:0] dcache_tlb_real_hits_lo =3'h0; 
    wire[2:0] dcache_tlb_real_hits_hi =3'h0; 
    wire[2:0] dcache_pma_checker_real_hits_lo =3'h0; 
    wire[2:0] dcache_pma_checker_real_hits_hi =3'h0; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_hi_lo_lo =3'h0; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_hi_lo_hi =3'h0; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_hi_hi_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_hi =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_hi =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_hi =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_lo =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_hi =3'h0; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_lo =3'h0; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_lo =3'h0; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_hi =3'h0; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_lo =3'h0; 
    wire[2:0] dcache_get_param =3'h0; 
    wire[2:0] dcache_put_opcode =3'h0; 
    wire[2:0] dcache_put_param =3'h0; 
    wire[2:0] dcache_putpartial_param =3'h0; 
    wire[2:0] dcache_atomics_a_1_param =3'h0; 
    wire[2:0] dcache_atomics_a_5_param =3'h0; 
    wire[17:0] dcache_dummyMeta_tag =18'h0; 
    wire[17:0] dcache_s2_meta_corrected_0_tag =18'h0; 
    wire[17:0] dcache_metaArb_io_in_1_bits_data_new_meta_tag =18'h0; 
    wire[17:0] dcache_metaArb_io_in_0_bits_data_meta_1_tag =18'h0; 
    wire[6:0] dcache_tlb_hr_array =7'h7F; 
    wire[6:0] dcache_tlb_hw_array =7'h7F; 
    wire[6:0] dcache_tlb_hx_array =7'h7F; 
    wire[6:0] dcache_pma_checker_hr_array =7'h7F; 
    wire[6:0] dcache_pma_checker_hw_array =7'h7F; 
    wire[6:0] dcache_pma_checker_hx_array =7'h7F; 
    wire[1:0] dcache_s2_victim_way =2'h1; 
    wire[1:0] dcache_dataArb_io_in_0_bits_wordMask_wordMask =2'h1; 
    wire[19:0] dcache_pma_checker_refill_ppn =20'h0; 
    wire[19:0] dcache_pma_checker_newEntry_ppn =20'h0; 
    wire[19:0] dcache_s1_meta_0 =20'h0; 
    wire[21:0] dcache_tlb_satp_ppn =22'h0; 
    wire[21:0] dcache_pma_checker_satp_ppn =22'h0; 
    wire[21:0] dcache_pma_checker_special_entry_data_0_hi_hi_hi =22'h0; 
    wire[21:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_hi =22'h0; 
    wire[21:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_hi =22'h0; 
    wire[21:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_hi =22'h0; 
    wire[21:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_hi =22'h0; 
    wire[21:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_hi =22'h0; 
    wire[7:0] dcache_flushCounterWrap =8'h1; 
    wire[8:0] dcache_flushCounterNext =9'h1; 
    wire[3:0] dcache_s0_req_mask =4'h0; 
    wire[3:0] dcache_nackResponseMessage_size =4'h0; 
    wire[3:0] dcache_cleanReleaseMessage_size =4'h0; 
    wire[3:0] dcache_dirtyReleaseMessage_size =4'h0; 
    wire[31:0] dcache_tl_out_c_bits_data =32'h0; 
    wire[31:0] dcache_s0_req_data =32'h0; 
    wire[31:0] dcache_get_data =32'h0; 
    wire[31:0] dcache_nackResponseMessage_address =32'h0; 
    wire[31:0] dcache_nackResponseMessage_data =32'h0; 
    wire[31:0] dcache_cleanReleaseMessage_address =32'h0; 
    wire[31:0] dcache_cleanReleaseMessage_data =32'h0; 
    wire[31:0] dcache_dirtyReleaseMessage_address =32'h0; 
    wire[31:0] dcache_dirtyReleaseMessage_data =32'h0; 
    wire[9:0] dcache_beats1_1 =10'h0; 
    wire[9:0] dcache_c_count =10'h0; 
    wire[9:0] dcache_io_cpu_perf_release_beats1 =10'h0; 
    wire[9:0] dcache_io_cpu_perf_release_count =10'h0; 
    wire[2:0] dcache_tl_out_c_bits_param =3'h5; 
    wire[2:0] dcache_nackResponseMessage_param =3'h5; 
    wire[2:0] dcache_dirtyReleaseMessage_opcode =3'h5; 
    wire[2:0] dcache_tl_out_c_bits_opcode =3'h4; 
    wire[2:0] dcache_get_opcode =3'h4; 
    wire[2:0] dcache_atomics_a_4_param =3'h4; 
    wire[2:0] dcache_nackResponseMessage_opcode =3'h4; 
    wire[2:0] dcache_cleanReleaseMessage_opcode =3'h4; 
    wire[2:0] dcache_atomics_a_opcode =3'h3; 
    wire[2:0] dcache_atomics_a_param =3'h3; 
    wire[2:0] dcache_atomics_a_1_opcode =3'h3; 
    wire[2:0] dcache_atomics_a_2_opcode =3'h3; 
    wire[2:0] dcache_atomics_a_3_opcode =3'h3; 
    wire[2:0] dcache_atomics_a_8_param =3'h3; 
    wire[2:0] dcache_atomics_a_3_param =3'h2; 
    wire[2:0] dcache_atomics_a_4_opcode =3'h2; 
    wire[2:0] dcache_atomics_a_5_opcode =3'h2; 
    wire[2:0] dcache_atomics_a_6_opcode =3'h2; 
    wire[2:0] dcache_atomics_a_7_opcode =3'h2; 
    wire[2:0] dcache_atomics_a_7_param =3'h2; 
    wire[2:0] dcache_atomics_a_8_opcode =3'h2; 
    wire[2:0] dcache_putpartial_opcode =3'h1; 
    wire[2:0] dcache_atomics_a_2_param =3'h1; 
    wire[2:0] dcache_atomics_a_6_param =3'h1; 
    wire[31:0] dcache_baseAddr =32'h80000000; 
    wire[5:0] dcache_tlb_stage2_bypass =6'h3F; 
    wire[5:0] dcache_tlb_gpa_hits_hit_mask =6'h3F; 
    wire[5:0] dcache_tlb_gpa_hits =6'h3F; 
    wire[5:0] dcache_pma_checker_stage2_bypass =6'h3F; 
    wire[5:0] dcache_pma_checker_gpa_hits_hit_mask =6'h3F; 
    wire[5:0] dcache_pma_checker_gpa_hits =6'h3F; 
    wire[6:0] dcache_tlb_lrscAllowed =7'h0; 
    wire[6:0] dcache_tlb_gf_ld_array =7'h0; 
    wire[6:0] dcache_tlb_gf_st_array =7'h0; 
    wire[6:0] dcache_tlb_gf_inst_array =7'h0; 
    wire[6:0] dcache_tlb_gpa_hits_need_gpa_mask =7'h0; 
    wire[6:0] dcache_pma_checker_lrscAllowed =7'h0; 
    wire[6:0] dcache_pma_checker_gf_ld_array =7'h0; 
    wire[6:0] dcache_pma_checker_gf_st_array =7'h0; 
    wire[6:0] dcache_pma_checker_gf_inst_array =7'h0; 
    wire[6:0] dcache_pma_checker_gpa_hits_need_gpa_mask =7'h0; 
    wire[30:0] dcache_pma_checker_special_entry_data_0_hi =31'h0; 
    wire[30:0] dcache_pma_checker_superpage_entries_0_data_0_hi =31'h0; 
    wire[30:0] dcache_pma_checker_superpage_entries_1_data_0_hi =31'h0; 
    wire[30:0] dcache_pma_checker_superpage_entries_2_data_0_hi =31'h0; 
    wire[30:0] dcache_pma_checker_superpage_entries_3_data_0_hi =31'h0; 
    wire[30:0] dcache_pma_checker_sectored_entries_0_0_data_hi =31'h0; 
    wire[20:0] dcache_pma_checker_special_entry_data_0_hi_hi_hi_hi =21'h0; 
    wire[20:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_hi_hi =21'h0; 
    wire[20:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_hi_hi =21'h0; 
    wire[20:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_hi_hi =21'h0; 
    wire[20:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_hi_hi =21'h0; 
    wire[20:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_hi_hi =21'h0; 
    wire[6:0] dcache_tlb_hits =7'h40; 
    wire[6:0] dcache_pma_checker_hits =7'h40; 
    wire dcache_nodeOut_a_deq_ready = dcache_nodeOut_a_ready ; 
    wire dcache_nodeOut_a_deq_valid ; 
    wire[2:0] dcache_nodeOut_a_deq_bits_opcode ; 
    wire[2:0] dcache_nodeOut_a_deq_bits_param ; 
    wire[3:0] dcache_nodeOut_a_deq_bits_size ; 
    wire[31:0] dcache_nodeOut_a_deq_bits_address ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_bufferable ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_modifiable ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_readalloc ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_writealloc ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_privileged ; 
    wire[3:0] dcache_nodeOut_a_deq_bits_mask ; 
    wire[31:0] dcache_nodeOut_a_deq_bits_data ; 
    wire dcache_e_sink = dcache_nodeOut_d_bits_sink ; 
    wire[31:0] dcache_s1_uncached_data_word = dcache_nodeOut_d_bits_data ; 
    wire[19:0] dcache_tlb_vpn = dcache_s1_tlb_req_vaddr [31:12]; 
    wire[19:0] dcache_tlb_ppn = dcache_tlb_vpn ; 
    wire dcache_tlb_priv_s = dcache_s1_tlb_req_prv [0]; 
    wire dcache_tlb_priv_uses_vm =~( dcache_s1_tlb_req_prv [1]); 
    wire[19:0] dcache_tlb_refill_ppn = dcache_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire[19:0] dcache_tlb_newEntry_ppn = dcache_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire[19:0] dcache_tlb_mpu_ppn = dcache_s1_tlb_req_vaddr [31:12]; 
    wire[11:0] dcache_tlb_io_resp_gpa_offset = dcache_s1_tlb_req_vaddr [11:0]; 
    wire[31:0] dcache_tlb_mpu_physaddr ={ dcache_tlb_mpu_ppn , dcache_tlb_io_resp_gpa_offset }; 
    wire[2:0] dcache_tlb_mpu_priv ={ dcache_io_ptw_status_debug , dcache_s1_tlb_req_prv }; 
    wire[19:0] dcache__GEN_0 ={ dcache_tlb_mpu_physaddr [31:14],~( dcache_tlb_mpu_physaddr [13:12])}; 
    wire[5:0] dcache__GEN_1 ={ dcache_tlb_mpu_physaddr [31:28],~( dcache_tlb_mpu_physaddr [27:26])}; 
    wire[9:0] dcache__GEN_2 = dcache_tlb_mpu_physaddr [25:16]^10'h200; 
    wire[15:0] dcache__GEN_3 ={ dcache_tlb_mpu_physaddr [31:26], dcache__GEN_2 }; 
    wire dcache__GEN_4 = dcache_tlb_mpu_physaddr [31:14]!=18'h20000; 
    wire[15:0] dcache__GEN_5 ={ dcache_tlb_mpu_physaddr [31:17],~( dcache_tlb_mpu_physaddr [16])}; 
    wire[2:0] dcache__GEN_6 ={ dcache_tlb_mpu_physaddr [31],~( dcache_tlb_mpu_physaddr [30:29])}; 
    wire dcache_tlb_legal_address =~(| dcache__GEN_0 )|~(| dcache__GEN_1 )|~(| dcache__GEN_3 )|~ dcache__GEN_4 |~(|( dcache_tlb_mpu_physaddr [31:12]))|~(| dcache__GEN_5 )|~(| dcache__GEN_6 ); 
    wire dcache_tlb_homogeneous =~(|( dcache_tlb_mpu_physaddr [31:12]))|~(| dcache__GEN_0 )|~(| dcache__GEN_5 )|~(| dcache__GEN_3 )|~(| dcache__GEN_1 )|~(| dcache__GEN_6 )|~ dcache__GEN_4 ; 
    wire dcache_tlb_deny_access_to_debug =~( dcache_tlb_mpu_priv [2])&~(|( dcache_tlb_mpu_physaddr [31:12])); 
    wire dcache_tlb_prot_r = dcache_tlb_legal_address &~ dcache_tlb_deny_access_to_debug & dcache__tlb_pmp_io_r ; 
    wire dcache_tlb_newEntry_pr = dcache_tlb_prot_r ; 
    wire[2:0] dcache__GEN_7 ={ dcache_tlb_mpu_physaddr [30], dcache_tlb_mpu_physaddr [27], dcache_tlb_mpu_physaddr [16]}; 
    wire[2:0] dcache__GEN_8 ={ dcache_tlb_mpu_physaddr [31:30],~( dcache_tlb_mpu_physaddr [27])}; 
    wire[1:0] dcache__GEN_9 ={ dcache_tlb_mpu_physaddr [31],~( dcache_tlb_mpu_physaddr [30])}; 
    wire dcache_tlb_prot_w = dcache_tlb_legal_address &(~(| dcache__GEN_7 )|~(| dcache__GEN_8 )|~(| dcache__GEN_9 ))&~ dcache_tlb_deny_access_to_debug & dcache__tlb_pmp_io_w ; 
    wire dcache_tlb_newEntry_pw = dcache_tlb_prot_w ; 
    wire dcache_tlb_prot_pp = dcache_tlb_legal_address &(~(| dcache__GEN_7 )|~(| dcache__GEN_8 )|~(| dcache__GEN_9 )); 
    wire dcache_tlb_newEntry_ppp = dcache_tlb_prot_pp ; 
    wire dcache_tlb_prot_al = dcache_tlb_legal_address &(~(| dcache__GEN_7 )|~(| dcache__GEN_8 )); 
    wire dcache_tlb_newEntry_pal = dcache_tlb_prot_al ; 
    wire dcache_tlb_prot_aa = dcache_tlb_legal_address &(~(| dcache__GEN_7 )|~(| dcache__GEN_8 )); 
    wire dcache_tlb_newEntry_paa = dcache_tlb_prot_aa ; 
    wire dcache_tlb_prot_x = dcache_tlb_legal_address &({ dcache_tlb_mpu_physaddr [30], dcache_tlb_mpu_physaddr [27], dcache_tlb_mpu_physaddr [25]}==3'h0|~(| dcache__GEN_9 ))&~ dcache_tlb_deny_access_to_debug & dcache__tlb_pmp_io_x ; 
    wire dcache_tlb_newEntry_px = dcache_tlb_prot_x ; 
    wire dcache_tlb_prot_eff = dcache_tlb_legal_address &({ dcache_tlb_mpu_physaddr [31:30], dcache_tlb_mpu_physaddr [27], dcache_tlb_mpu_physaddr [25], dcache_tlb_mpu_physaddr [16], dcache_tlb_mpu_physaddr [13]}==6'h0|{ dcache_tlb_mpu_physaddr [31:30], dcache_tlb_mpu_physaddr [27], dcache__GEN_2 [9], dcache_tlb_mpu_physaddr [16]}==5'h0|~(| dcache__GEN_8 )|~(| dcache__GEN_9 )); 
    wire dcache_tlb_newEntry_eff = dcache_tlb_prot_eff ; 
    wire[1:0] dcache_tlb_hitsVec_idx = dcache_tlb_vpn [1:0]; 
    wire dcache_tlb_newEntry_g = dcache_io_ptw_resp_bits_pte_g & dcache_io_ptw_resp_bits_pte_v ; 
    wire dcache_tlb_newEntry_sr = dcache_io_ptw_resp_bits_pte_v &( dcache_io_ptw_resp_bits_pte_r | dcache_io_ptw_resp_bits_pte_x &~ dcache_io_ptw_resp_bits_pte_w )& dcache_io_ptw_resp_bits_pte_a & dcache_io_ptw_resp_bits_pte_r ; 
    wire dcache_tlb_newEntry_sw = dcache_io_ptw_resp_bits_pte_v &( dcache_io_ptw_resp_bits_pte_r | dcache_io_ptw_resp_bits_pte_x &~ dcache_io_ptw_resp_bits_pte_w )& dcache_io_ptw_resp_bits_pte_a & dcache_io_ptw_resp_bits_pte_w & dcache_io_ptw_resp_bits_pte_d ; 
    wire dcache_tlb_newEntry_sx = dcache_io_ptw_resp_bits_pte_v &( dcache_io_ptw_resp_bits_pte_r | dcache_io_ptw_resp_bits_pte_x &~ dcache_io_ptw_resp_bits_pte_w )& dcache_io_ptw_resp_bits_pte_a & dcache_io_ptw_resp_bits_pte_x ; 
    wire[1:0] dcache__GEN_10 ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_lo_hi_hi ; 
  assign  dcache_tlb_special_entry_data_0_lo_lo_hi_hi = dcache__GEN_10 ; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_lo_lo_hi_hi = dcache__GEN_10 ; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_lo_lo_hi_hi = dcache__GEN_10 ; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_lo_lo_hi_hi = dcache__GEN_10 ; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_lo_lo_hi_hi = dcache__GEN_10 ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_lo_hi_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_lo_lo_hi_hi = dcache__GEN_10 ; 
    wire[2:0] dcache_tlb_special_entry_data_0_lo_lo_hi ={ dcache_tlb_special_entry_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_special_entry_data_0_lo_lo ={ dcache_tlb_special_entry_data_0_lo_lo_hi ,2'h0}; 
    wire[1:0] dcache__GEN_11 ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_hi_lo_hi ; 
  assign  dcache_tlb_special_entry_data_0_lo_hi_lo_hi = dcache__GEN_11 ; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_lo_hi_lo_hi = dcache__GEN_11 ; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_lo_hi_lo_hi = dcache__GEN_11 ; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_lo_hi_lo_hi = dcache__GEN_11 ; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_lo_hi_lo_hi = dcache__GEN_11 ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_lo_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_lo_hi_lo_hi = dcache__GEN_11 ; 
    wire[2:0] dcache_tlb_special_entry_data_0_lo_hi_lo ={ dcache_tlb_special_entry_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache__GEN_12 ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_hi_hi_hi ; 
  assign  dcache_tlb_special_entry_data_0_lo_hi_hi_hi = dcache__GEN_12 ; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_lo_hi_hi_hi = dcache__GEN_12 ; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_lo_hi_hi_hi = dcache__GEN_12 ; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_lo_hi_hi_hi = dcache__GEN_12 ; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_lo_hi_hi_hi = dcache__GEN_12 ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_hi_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_lo_hi_hi_hi = dcache__GEN_12 ; 
    wire[2:0] dcache_tlb_special_entry_data_0_lo_hi_hi ={ dcache_tlb_special_entry_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_special_entry_data_0_lo_hi ={ dcache_tlb_special_entry_data_0_lo_hi_hi , dcache_tlb_special_entry_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_special_entry_data_0_lo ={ dcache_tlb_special_entry_data_0_lo_hi , dcache_tlb_special_entry_data_0_lo_lo }; 
    wire[1:0] dcache__GEN_13 ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[1:0] dcache_tlb_special_entry_data_0_hi_lo_lo_hi ; 
  assign  dcache_tlb_special_entry_data_0_hi_lo_lo_hi = dcache__GEN_13 ; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_lo_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_hi_lo_lo_hi = dcache__GEN_13 ; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_lo_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_hi_lo_lo_hi = dcache__GEN_13 ; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_lo_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_hi_lo_lo_hi = dcache__GEN_13 ; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_lo_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_hi_lo_lo_hi = dcache__GEN_13 ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_lo_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_hi_lo_lo_hi = dcache__GEN_13 ; 
    wire[2:0] dcache_tlb_special_entry_data_0_hi_lo_lo ={ dcache_tlb_special_entry_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache__GEN_14 ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[1:0] dcache_tlb_special_entry_data_0_hi_lo_hi_hi ; 
  assign  dcache_tlb_special_entry_data_0_hi_lo_hi_hi = dcache__GEN_14 ; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_hi_lo_hi_hi = dcache__GEN_14 ; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_hi_lo_hi_hi = dcache__GEN_14 ; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_hi_lo_hi_hi = dcache__GEN_14 ; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_hi_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_hi_lo_hi_hi = dcache__GEN_14 ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_hi_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_hi_lo_hi_hi = dcache__GEN_14 ; 
    wire[2:0] dcache_tlb_special_entry_data_0_hi_lo_hi ={ dcache_tlb_special_entry_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_special_entry_data_0_hi_lo ={ dcache_tlb_special_entry_data_0_hi_lo_hi , dcache_tlb_special_entry_data_0_hi_lo_lo }; 
    wire[1:0] dcache__GEN_15 ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[1:0] dcache_tlb_special_entry_data_0_hi_hi_lo_hi ; 
  assign  dcache_tlb_special_entry_data_0_hi_hi_lo_hi = dcache__GEN_15 ; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_hi_hi_lo_hi = dcache__GEN_15 ; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_hi_hi_lo_hi = dcache__GEN_15 ; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_hi_hi_lo_hi = dcache__GEN_15 ; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_lo_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_hi_hi_lo_hi = dcache__GEN_15 ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_lo_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_hi_hi_lo_hi = dcache__GEN_15 ; 
    wire[2:0] dcache_tlb_special_entry_data_0_hi_hi_lo ={ dcache_tlb_special_entry_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache__GEN_16 ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[20:0] dcache_tlb_special_entry_data_0_hi_hi_hi_hi ; 
  assign  dcache_tlb_special_entry_data_0_hi_hi_hi_hi = dcache__GEN_16 ; 
    wire[20:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_0_data_0_hi_hi_hi_hi = dcache__GEN_16 ; 
    wire[20:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_1_data_0_hi_hi_hi_hi = dcache__GEN_16 ; 
    wire[20:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_2_data_0_hi_hi_hi_hi = dcache__GEN_16 ; 
    wire[20:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_hi_hi ; 
  assign  dcache_tlb_superpage_entries_3_data_0_hi_hi_hi_hi = dcache__GEN_16 ; 
    wire[20:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_hi_hi ; 
  assign  dcache_tlb_sectored_entries_0_0_data_hi_hi_hi_hi = dcache__GEN_16 ; 
    wire[21:0] dcache_tlb_special_entry_data_0_hi_hi_hi ={ dcache_tlb_special_entry_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_special_entry_data_0_hi_hi ={ dcache_tlb_special_entry_data_0_hi_hi_hi , dcache_tlb_special_entry_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_special_entry_data_0_hi ={ dcache_tlb_special_entry_data_0_hi_hi , dcache_tlb_special_entry_data_0_hi_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_0_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_0_data_0_lo_lo ={ dcache_tlb_superpage_entries_0_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_0_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_0_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_0_data_0_lo_hi ={ dcache_tlb_superpage_entries_0_data_0_lo_hi_hi , dcache_tlb_superpage_entries_0_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_0_data_0_lo ={ dcache_tlb_superpage_entries_0_data_0_lo_hi , dcache_tlb_superpage_entries_0_data_0_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_0_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_0_data_0_hi_lo ={ dcache_tlb_superpage_entries_0_data_0_hi_lo_hi , dcache_tlb_superpage_entries_0_data_0_hi_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_0_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[21:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_0_data_0_hi_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_hi_hi , dcache_tlb_superpage_entries_0_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_0_data_0_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_hi , dcache_tlb_superpage_entries_0_data_0_hi_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_1_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_1_data_0_lo_lo ={ dcache_tlb_superpage_entries_1_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_1_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_1_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_1_data_0_lo_hi ={ dcache_tlb_superpage_entries_1_data_0_lo_hi_hi , dcache_tlb_superpage_entries_1_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_1_data_0_lo ={ dcache_tlb_superpage_entries_1_data_0_lo_hi , dcache_tlb_superpage_entries_1_data_0_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_1_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_1_data_0_hi_lo ={ dcache_tlb_superpage_entries_1_data_0_hi_lo_hi , dcache_tlb_superpage_entries_1_data_0_hi_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_1_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[21:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_1_data_0_hi_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_hi_hi , dcache_tlb_superpage_entries_1_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_1_data_0_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_hi , dcache_tlb_superpage_entries_1_data_0_hi_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_2_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_2_data_0_lo_lo ={ dcache_tlb_superpage_entries_2_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_2_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_2_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_2_data_0_lo_hi ={ dcache_tlb_superpage_entries_2_data_0_lo_hi_hi , dcache_tlb_superpage_entries_2_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_2_data_0_lo ={ dcache_tlb_superpage_entries_2_data_0_lo_hi , dcache_tlb_superpage_entries_2_data_0_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_2_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_2_data_0_hi_lo ={ dcache_tlb_superpage_entries_2_data_0_hi_lo_hi , dcache_tlb_superpage_entries_2_data_0_hi_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_2_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[21:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_2_data_0_hi_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_hi_hi , dcache_tlb_superpage_entries_2_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_2_data_0_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_hi , dcache_tlb_superpage_entries_2_data_0_hi_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_3_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_3_data_0_lo_lo ={ dcache_tlb_superpage_entries_3_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_3_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_3_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_3_data_0_lo_hi ={ dcache_tlb_superpage_entries_3_data_0_lo_hi_hi , dcache_tlb_superpage_entries_3_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_3_data_0_lo ={ dcache_tlb_superpage_entries_3_data_0_lo_hi , dcache_tlb_superpage_entries_3_data_0_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_3_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_3_data_0_hi_lo ={ dcache_tlb_superpage_entries_3_data_0_hi_lo_hi , dcache_tlb_superpage_entries_3_data_0_hi_lo_lo }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_3_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[21:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_3_data_0_hi_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_hi_hi , dcache_tlb_superpage_entries_3_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_3_data_0_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_hi , dcache_tlb_superpage_entries_3_data_0_hi_lo }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_lo_lo_hi ={ dcache_tlb_sectored_entries_0_0_data_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_sectored_entries_0_0_data_lo_lo ={ dcache_tlb_sectored_entries_0_0_data_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_lo ={ dcache_tlb_sectored_entries_0_0_data_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_hi ={ dcache_tlb_sectored_entries_0_0_data_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_sectored_entries_0_0_data_lo_hi ={ dcache_tlb_sectored_entries_0_0_data_lo_hi_hi , dcache_tlb_sectored_entries_0_0_data_lo_hi_lo }; 
    wire[10:0] dcache_tlb_sectored_entries_0_0_data_lo ={ dcache_tlb_sectored_entries_0_0_data_lo_hi , dcache_tlb_sectored_entries_0_0_data_lo_lo }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_lo ={ dcache_tlb_sectored_entries_0_0_data_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_sectored_entries_0_0_data_hi_lo ={ dcache_tlb_sectored_entries_0_0_data_hi_lo_hi , dcache_tlb_sectored_entries_0_0_data_hi_lo_lo }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_lo ={ dcache_tlb_sectored_entries_0_0_data_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[21:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_sectored_entries_0_0_data_hi_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_hi_hi , dcache_tlb_sectored_entries_0_0_data_hi_hi_lo }; 
    wire[30:0] dcache_tlb_sectored_entries_0_0_data_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_hi , dcache_tlb_sectored_entries_0_0_data_hi_lo }; 
    wire[1:0] dcache_tlb_ptw_ae_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_ae_ptw , dcache__tlb_entries_barrier_1_io_y_ae_ptw }; 
    wire[2:0] dcache_tlb_ptw_ae_array_lo ={ dcache_tlb_ptw_ae_array_lo_hi , dcache__tlb_entries_barrier_io_y_ae_ptw }; 
    wire[1:0] dcache_tlb_ptw_ae_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_ae_ptw , dcache__tlb_entries_barrier_4_io_y_ae_ptw }; 
    wire[2:0] dcache_tlb_ptw_ae_array_hi ={ dcache_tlb_ptw_ae_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_ae_ptw }; 
    wire[6:0] dcache_tlb_ptw_ae_array ={1'h0, dcache_tlb_ptw_ae_array_hi , dcache_tlb_ptw_ae_array_lo }; 
    wire[1:0] dcache_tlb_final_ae_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_ae_final , dcache__tlb_entries_barrier_1_io_y_ae_final }; 
    wire[2:0] dcache_tlb_final_ae_array_lo ={ dcache_tlb_final_ae_array_lo_hi , dcache__tlb_entries_barrier_io_y_ae_final }; 
    wire[1:0] dcache_tlb_final_ae_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_ae_final , dcache__tlb_entries_barrier_4_io_y_ae_final }; 
    wire[2:0] dcache_tlb_final_ae_array_hi ={ dcache_tlb_final_ae_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_ae_final }; 
    wire[6:0] dcache_tlb_final_ae_array ={1'h0, dcache_tlb_final_ae_array_hi , dcache_tlb_final_ae_array_lo }; 
    wire[1:0] dcache_tlb_ptw_pf_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_pf , dcache__tlb_entries_barrier_1_io_y_pf }; 
    wire[2:0] dcache_tlb_ptw_pf_array_lo ={ dcache_tlb_ptw_pf_array_lo_hi , dcache__tlb_entries_barrier_io_y_pf }; 
    wire[1:0] dcache_tlb_ptw_pf_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_pf , dcache__tlb_entries_barrier_4_io_y_pf }; 
    wire[2:0] dcache_tlb_ptw_pf_array_hi ={ dcache_tlb_ptw_pf_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_pf }; 
    wire[6:0] dcache_tlb_ptw_pf_array ={1'h0, dcache_tlb_ptw_pf_array_hi , dcache_tlb_ptw_pf_array_lo }; 
    wire[1:0] dcache_tlb_ptw_gf_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_gf , dcache__tlb_entries_barrier_1_io_y_gf }; 
    wire[2:0] dcache_tlb_ptw_gf_array_lo ={ dcache_tlb_ptw_gf_array_lo_hi , dcache__tlb_entries_barrier_io_y_gf }; 
    wire[1:0] dcache_tlb_ptw_gf_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_gf , dcache__tlb_entries_barrier_4_io_y_gf }; 
    wire[2:0] dcache_tlb_ptw_gf_array_hi ={ dcache_tlb_ptw_gf_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_gf }; 
    wire[6:0] dcache_tlb_ptw_gf_array ={1'h0, dcache_tlb_ptw_gf_array_hi , dcache_tlb_ptw_gf_array_lo }; 
    wire[1:0] dcache__GEN_17 ={ dcache__tlb_entries_barrier_2_io_y_u , dcache__tlb_entries_barrier_1_io_y_u }; 
    wire[1:0] dcache_tlb_priv_rw_ok_lo_hi ; 
  assign  dcache_tlb_priv_rw_ok_lo_hi = dcache__GEN_17 ; 
    wire[1:0] dcache_tlb_priv_rw_ok_lo_hi_1 ; 
  assign  dcache_tlb_priv_rw_ok_lo_hi_1 = dcache__GEN_17 ; 
    wire[1:0] dcache_tlb_priv_x_ok_lo_hi ; 
  assign  dcache_tlb_priv_x_ok_lo_hi = dcache__GEN_17 ; 
    wire[1:0] dcache_tlb_priv_x_ok_lo_hi_1 ; 
  assign  dcache_tlb_priv_x_ok_lo_hi_1 = dcache__GEN_17 ; 
    wire[2:0] dcache_tlb_priv_rw_ok_lo ={ dcache_tlb_priv_rw_ok_lo_hi , dcache__tlb_entries_barrier_io_y_u }; 
    wire[1:0] dcache__GEN_18 ={ dcache__tlb_entries_barrier_5_io_y_u , dcache__tlb_entries_barrier_4_io_y_u }; 
    wire[1:0] dcache_tlb_priv_rw_ok_hi_hi ; 
  assign  dcache_tlb_priv_rw_ok_hi_hi = dcache__GEN_18 ; 
    wire[1:0] dcache_tlb_priv_rw_ok_hi_hi_1 ; 
  assign  dcache_tlb_priv_rw_ok_hi_hi_1 = dcache__GEN_18 ; 
    wire[1:0] dcache_tlb_priv_x_ok_hi_hi ; 
  assign  dcache_tlb_priv_x_ok_hi_hi = dcache__GEN_18 ; 
    wire[1:0] dcache_tlb_priv_x_ok_hi_hi_1 ; 
  assign  dcache_tlb_priv_x_ok_hi_hi_1 = dcache__GEN_18 ; 
    wire[2:0] dcache_tlb_priv_rw_ok_hi ={ dcache_tlb_priv_rw_ok_hi_hi , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[2:0] dcache_tlb_priv_rw_ok_lo_1 ={ dcache_tlb_priv_rw_ok_lo_hi_1 , dcache__tlb_entries_barrier_io_y_u }; 
    wire[2:0] dcache_tlb_priv_rw_ok_hi_1 ={ dcache_tlb_priv_rw_ok_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_tlb_priv_rw_ok =( dcache_tlb_priv_s  ? 6'h0:{ dcache_tlb_priv_rw_ok_hi , dcache_tlb_priv_rw_ok_lo })|( dcache_tlb_priv_s  ? ~{ dcache_tlb_priv_rw_ok_hi_1 , dcache_tlb_priv_rw_ok_lo_1 }:6'h0); 
    wire[2:0] dcache_tlb_priv_x_ok_lo ={ dcache_tlb_priv_x_ok_lo_hi , dcache__tlb_entries_barrier_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_hi ={ dcache_tlb_priv_x_ok_hi_hi , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_lo_1 ={ dcache_tlb_priv_x_ok_lo_hi_1 , dcache__tlb_entries_barrier_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_hi_1 ={ dcache_tlb_priv_x_ok_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_tlb_priv_x_ok = dcache_tlb_priv_s  ? ~{ dcache_tlb_priv_x_ok_hi , dcache_tlb_priv_x_ok_lo }:{ dcache_tlb_priv_x_ok_hi_1 , dcache_tlb_priv_x_ok_lo_1 }; 
    wire[1:0] dcache_tlb_stage1_bypass_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_ae_stage2 , dcache__tlb_entries_barrier_1_io_y_ae_stage2 }; 
    wire[2:0] dcache_tlb_stage1_bypass_lo ={ dcache_tlb_stage1_bypass_lo_hi , dcache__tlb_entries_barrier_io_y_ae_stage2 }; 
    wire[1:0] dcache_tlb_stage1_bypass_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_ae_stage2 , dcache__tlb_entries_barrier_4_io_y_ae_stage2 }; 
    wire[2:0] dcache_tlb_stage1_bypass_hi ={ dcache_tlb_stage1_bypass_hi_hi , dcache__tlb_entries_barrier_3_io_y_ae_stage2 }; 
    wire[1:0] dcache_tlb_r_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_sr , dcache__tlb_entries_barrier_1_io_y_sr }; 
    wire[2:0] dcache_tlb_r_array_lo ={ dcache_tlb_r_array_lo_hi , dcache__tlb_entries_barrier_io_y_sr }; 
    wire[1:0] dcache_tlb_r_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_sr , dcache__tlb_entries_barrier_4_io_y_sr }; 
    wire[2:0] dcache_tlb_r_array_hi ={ dcache_tlb_r_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_sr }; 
    wire[1:0] dcache__GEN_19 ={ dcache__tlb_entries_barrier_2_io_y_sx , dcache__tlb_entries_barrier_1_io_y_sx }; 
    wire[1:0] dcache_tlb_r_array_lo_hi_1 ; 
  assign  dcache_tlb_r_array_lo_hi_1 = dcache__GEN_19 ; 
    wire[1:0] dcache_tlb_x_array_lo_hi ; 
  assign  dcache_tlb_x_array_lo_hi = dcache__GEN_19 ; 
    wire[2:0] dcache_tlb_r_array_lo_1 ={ dcache_tlb_r_array_lo_hi_1 , dcache__tlb_entries_barrier_io_y_sx }; 
    wire[1:0] dcache__GEN_20 ={ dcache__tlb_entries_barrier_5_io_y_sx , dcache__tlb_entries_barrier_4_io_y_sx }; 
    wire[1:0] dcache_tlb_r_array_hi_hi_1 ; 
  assign  dcache_tlb_r_array_hi_hi_1 = dcache__GEN_20 ; 
    wire[1:0] dcache_tlb_x_array_hi_hi ; 
  assign  dcache_tlb_x_array_hi_hi = dcache__GEN_20 ; 
    wire[2:0] dcache_tlb_r_array_hi_1 ={ dcache_tlb_r_array_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_tlb_r_array ={1'h1, dcache_tlb_priv_rw_ok &{ dcache_tlb_r_array_hi , dcache_tlb_r_array_lo }}; 
    wire[1:0] dcache_tlb_w_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_sw , dcache__tlb_entries_barrier_1_io_y_sw }; 
    wire[2:0] dcache_tlb_w_array_lo ={ dcache_tlb_w_array_lo_hi , dcache__tlb_entries_barrier_io_y_sw }; 
    wire[1:0] dcache_tlb_w_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_sw , dcache__tlb_entries_barrier_4_io_y_sw }; 
    wire[2:0] dcache_tlb_w_array_hi ={ dcache_tlb_w_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_sw }; 
    wire[6:0] dcache_tlb_w_array ={1'h1, dcache_tlb_priv_rw_ok &{ dcache_tlb_w_array_hi , dcache_tlb_w_array_lo }}; 
    wire[2:0] dcache_tlb_x_array_lo ={ dcache_tlb_x_array_lo_hi , dcache__tlb_entries_barrier_io_y_sx }; 
    wire[2:0] dcache_tlb_x_array_hi ={ dcache_tlb_x_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_tlb_x_array ={1'h1, dcache_tlb_priv_x_ok &{ dcache_tlb_x_array_hi , dcache_tlb_x_array_lo }}; 
    wire[1:0] dcache_tlb_hr_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_hr , dcache__tlb_entries_barrier_1_io_y_hr }; 
    wire[2:0] dcache_tlb_hr_array_lo ={ dcache_tlb_hr_array_lo_hi , dcache__tlb_entries_barrier_io_y_hr }; 
    wire[1:0] dcache_tlb_hr_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_hr , dcache__tlb_entries_barrier_4_io_y_hr }; 
    wire[2:0] dcache_tlb_hr_array_hi ={ dcache_tlb_hr_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_hr }; 
    wire[1:0] dcache__GEN_21 ={ dcache__tlb_entries_barrier_2_io_y_hx , dcache__tlb_entries_barrier_1_io_y_hx }; 
    wire[1:0] dcache_tlb_hr_array_lo_hi_1 ; 
  assign  dcache_tlb_hr_array_lo_hi_1 = dcache__GEN_21 ; 
    wire[1:0] dcache_tlb_hx_array_lo_hi ; 
  assign  dcache_tlb_hx_array_lo_hi = dcache__GEN_21 ; 
    wire[2:0] dcache_tlb_hr_array_lo_1 ={ dcache_tlb_hr_array_lo_hi_1 , dcache__tlb_entries_barrier_io_y_hx }; 
    wire[1:0] dcache__GEN_22 ={ dcache__tlb_entries_barrier_5_io_y_hx , dcache__tlb_entries_barrier_4_io_y_hx }; 
    wire[1:0] dcache_tlb_hr_array_hi_hi_1 ; 
  assign  dcache_tlb_hr_array_hi_hi_1 = dcache__GEN_22 ; 
    wire[1:0] dcache_tlb_hx_array_hi_hi ; 
  assign  dcache_tlb_hx_array_hi_hi = dcache__GEN_22 ; 
    wire[2:0] dcache_tlb_hr_array_hi_1 ={ dcache_tlb_hr_array_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_hx }; 
    wire[1:0] dcache_tlb_hw_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_hw , dcache__tlb_entries_barrier_1_io_y_hw }; 
    wire[2:0] dcache_tlb_hw_array_lo ={ dcache_tlb_hw_array_lo_hi , dcache__tlb_entries_barrier_io_y_hw }; 
    wire[1:0] dcache_tlb_hw_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_hw , dcache__tlb_entries_barrier_4_io_y_hw }; 
    wire[2:0] dcache_tlb_hw_array_hi ={ dcache_tlb_hw_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_hw }; 
    wire[2:0] dcache_tlb_hx_array_lo ={ dcache_tlb_hx_array_lo_hi , dcache__tlb_entries_barrier_io_y_hx }; 
    wire[2:0] dcache_tlb_hx_array_hi ={ dcache_tlb_hx_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_hx }; 
    wire[1:0] dcache_tlb_pr_array_lo ={ dcache__tlb_entries_barrier_1_io_y_pr , dcache__tlb_entries_barrier_io_y_pr }; 
    wire[1:0] dcache_tlb_pr_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_pr , dcache__tlb_entries_barrier_3_io_y_pr }; 
    wire[2:0] dcache_tlb_pr_array_hi ={ dcache_tlb_pr_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_pr }; 
    wire[6:0] dcache_tlb__pr_array_T_4 = dcache_tlb_ptw_ae_array | dcache_tlb_final_ae_array ; 
    wire[6:0] dcache_tlb_pr_array ={{2{ dcache_tlb_prot_r }}, dcache_tlb_pr_array_hi , dcache_tlb_pr_array_lo }&~ dcache_tlb__pr_array_T_4 ; 
    wire[1:0] dcache_tlb_pw_array_lo ={ dcache__tlb_entries_barrier_1_io_y_pw , dcache__tlb_entries_barrier_io_y_pw }; 
    wire[1:0] dcache_tlb_pw_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_pw , dcache__tlb_entries_barrier_3_io_y_pw }; 
    wire[2:0] dcache_tlb_pw_array_hi ={ dcache_tlb_pw_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_pw }; 
    wire[6:0] dcache_tlb_pw_array ={{2{ dcache_tlb_prot_w }}, dcache_tlb_pw_array_hi , dcache_tlb_pw_array_lo }&~ dcache_tlb__pr_array_T_4 ; 
    wire[1:0] dcache_tlb_px_array_lo ={ dcache__tlb_entries_barrier_1_io_y_px , dcache__tlb_entries_barrier_io_y_px }; 
    wire[1:0] dcache_tlb_px_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_px , dcache__tlb_entries_barrier_3_io_y_px }; 
    wire[2:0] dcache_tlb_px_array_hi ={ dcache_tlb_px_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_px }; 
    wire[6:0] dcache_tlb_px_array ={{2{ dcache_tlb_prot_x }}, dcache_tlb_px_array_hi , dcache_tlb_px_array_lo }&~ dcache_tlb__pr_array_T_4 ; 
    wire[1:0] dcache_tlb_eff_array_lo ={ dcache__tlb_entries_barrier_1_io_y_eff , dcache__tlb_entries_barrier_io_y_eff }; 
    wire[1:0] dcache_tlb_eff_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_eff , dcache__tlb_entries_barrier_3_io_y_eff }; 
    wire[2:0] dcache_tlb_eff_array_hi ={ dcache_tlb_eff_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_eff }; 
    wire[6:0] dcache_tlb_eff_array ={{2{ dcache_tlb_prot_eff }}, dcache_tlb_eff_array_hi , dcache_tlb_eff_array_lo }; 
    wire[1:0] dcache__GEN_23 ={ dcache__tlb_entries_barrier_1_io_y_c , dcache__tlb_entries_barrier_io_y_c }; 
    wire[1:0] dcache_tlb_c_array_lo ; 
  assign  dcache_tlb_c_array_lo = dcache__GEN_23 ; 
    wire[1:0] dcache_tlb_prefetchable_array_lo ; 
  assign  dcache_tlb_prefetchable_array_lo = dcache__GEN_23 ; 
    wire[1:0] dcache__GEN_24 ={ dcache__tlb_entries_barrier_4_io_y_c , dcache__tlb_entries_barrier_3_io_y_c }; 
    wire[1:0] dcache_tlb_c_array_hi_hi ; 
  assign  dcache_tlb_c_array_hi_hi = dcache__GEN_24 ; 
    wire[1:0] dcache_tlb_prefetchable_array_hi_hi ; 
  assign  dcache_tlb_prefetchable_array_hi_hi = dcache__GEN_24 ; 
    wire[2:0] dcache_tlb_c_array_hi ={ dcache_tlb_c_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_tlb_c_array ={2'h0, dcache_tlb_c_array_hi , dcache_tlb_c_array_lo }; 
    wire[1:0] dcache_tlb_ppp_array_lo ={ dcache__tlb_entries_barrier_1_io_y_ppp , dcache__tlb_entries_barrier_io_y_ppp }; 
    wire[1:0] dcache_tlb_ppp_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_ppp , dcache__tlb_entries_barrier_3_io_y_ppp }; 
    wire[2:0] dcache_tlb_ppp_array_hi ={ dcache_tlb_ppp_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_ppp }; 
    wire[6:0] dcache_tlb_ppp_array ={{2{ dcache_tlb_prot_pp }}, dcache_tlb_ppp_array_hi , dcache_tlb_ppp_array_lo }; 
    wire[1:0] dcache_tlb_paa_array_lo ={ dcache__tlb_entries_barrier_1_io_y_paa , dcache__tlb_entries_barrier_io_y_paa }; 
    wire[1:0] dcache_tlb_paa_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_paa , dcache__tlb_entries_barrier_3_io_y_paa }; 
    wire[2:0] dcache_tlb_paa_array_hi ={ dcache_tlb_paa_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_paa }; 
    wire[6:0] dcache_tlb_paa_array ={{2{ dcache_tlb_prot_aa }}, dcache_tlb_paa_array_hi , dcache_tlb_paa_array_lo }; 
    wire[1:0] dcache_tlb_pal_array_lo ={ dcache__tlb_entries_barrier_1_io_y_pal , dcache__tlb_entries_barrier_io_y_pal }; 
    wire[1:0] dcache_tlb_pal_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_pal , dcache__tlb_entries_barrier_3_io_y_pal }; 
    wire[2:0] dcache_tlb_pal_array_hi ={ dcache_tlb_pal_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_pal }; 
    wire[6:0] dcache_tlb_pal_array ={{2{ dcache_tlb_prot_al }}, dcache_tlb_pal_array_hi , dcache_tlb_pal_array_lo }; 
    wire[6:0] dcache_tlb_ppp_array_if_cached = dcache_tlb_ppp_array | dcache_tlb_c_array ; 
    wire[6:0] dcache_tlb_paa_array_if_cached = dcache_tlb_paa_array | dcache_tlb_c_array ; 
    wire[6:0] dcache_tlb_pal_array_if_cached = dcache_tlb_pal_array | dcache_tlb_c_array ; 
    wire[2:0] dcache_tlb_prefetchable_array_hi ={ dcache_tlb_prefetchable_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_tlb_prefetchable_array ={2'h0, dcache_tlb_prefetchable_array_hi , dcache_tlb_prefetchable_array_lo }; 
    wire dcache_tlb_misaligned =|( dcache_s1_tlb_req_vaddr [3:0]&(4'h1<< dcache_s1_tlb_req_size )-4'h1); 
    wire dcache_tlb__cmd_lrsc_T = dcache_s1_tlb_req_cmd ==5'h6; 
    wire dcache_tlb__cmd_lrsc_T_1 = dcache_s1_tlb_req_cmd ==5'h7; 
    wire dcache_tlb_cmd_lrsc = dcache_tlb__cmd_lrsc_T | dcache_tlb__cmd_lrsc_T_1 ; 
    wire dcache_tlb__cmd_read_T_7 = dcache_s1_tlb_req_cmd ==5'h4; 
    wire dcache_tlb__cmd_read_T_8 = dcache_s1_tlb_req_cmd ==5'h9; 
    wire dcache_tlb__cmd_read_T_9 = dcache_s1_tlb_req_cmd ==5'hA; 
    wire dcache_tlb__cmd_read_T_10 = dcache_s1_tlb_req_cmd ==5'hB; 
    wire dcache_tlb_cmd_amo_logical = dcache_tlb__cmd_read_T_7 | dcache_tlb__cmd_read_T_8 | dcache_tlb__cmd_read_T_9 | dcache_tlb__cmd_read_T_10 ; 
    wire dcache_tlb__cmd_read_T_14 = dcache_s1_tlb_req_cmd ==5'h8; 
    wire dcache_tlb__cmd_read_T_15 = dcache_s1_tlb_req_cmd ==5'hC; 
    wire dcache_tlb__cmd_read_T_16 = dcache_s1_tlb_req_cmd ==5'hD; 
    wire dcache_tlb__cmd_read_T_17 = dcache_s1_tlb_req_cmd ==5'hE; 
    wire dcache_tlb__cmd_read_T_18 = dcache_s1_tlb_req_cmd ==5'hF; 
    wire dcache_tlb_cmd_amo_arithmetic = dcache_tlb__cmd_read_T_14 | dcache_tlb__cmd_read_T_15 | dcache_tlb__cmd_read_T_16 | dcache_tlb__cmd_read_T_17 | dcache_tlb__cmd_read_T_18 ; 
    wire dcache_tlb_cmd_put_partial = dcache_s1_tlb_req_cmd ==5'h11; 
    wire dcache_tlb_cmd_read = dcache_s1_tlb_req_cmd ==5'h0| dcache_s1_tlb_req_cmd ==5'h10| dcache_tlb__cmd_lrsc_T | dcache_tlb__cmd_lrsc_T_1 | dcache_tlb__cmd_read_T_7 | dcache_tlb__cmd_read_T_8 | dcache_tlb__cmd_read_T_9 | dcache_tlb__cmd_read_T_10 | dcache_tlb__cmd_read_T_14 | dcache_tlb__cmd_read_T_15 | dcache_tlb__cmd_read_T_16 | dcache_tlb__cmd_read_T_17 | dcache_tlb__cmd_read_T_18 ; 
    wire dcache_tlb_cmd_write = dcache_s1_tlb_req_cmd ==5'h1| dcache_tlb_cmd_put_partial | dcache_tlb__cmd_lrsc_T_1 | dcache_tlb__cmd_read_T_7 | dcache_tlb__cmd_read_T_8 | dcache_tlb__cmd_read_T_9 | dcache_tlb__cmd_read_T_10 | dcache_tlb__cmd_read_T_14 | dcache_tlb__cmd_read_T_15 | dcache_tlb__cmd_read_T_16 | dcache_tlb__cmd_read_T_17 | dcache_tlb__cmd_read_T_18 ; 
    wire dcache_tlb_cmd_write_perms = dcache_tlb_cmd_write | dcache_s1_tlb_req_cmd ==5'h5| dcache_s1_tlb_req_cmd ==5'h17; 
    wire[6:0] dcache_tlb_ae_array =( dcache_tlb_misaligned  ?  dcache_tlb_eff_array :7'h0)|{7{ dcache_tlb_cmd_lrsc }}; 
    wire[6:0] dcache_tlb_ae_ld_array = dcache_tlb_cmd_read  ?  dcache_tlb_ae_array |~ dcache_tlb_pr_array :7'h0; 
    wire[6:0] dcache_tlb_ae_st_array =( dcache_tlb_cmd_write_perms  ?  dcache_tlb_ae_array |~ dcache_tlb_pw_array :7'h0)|( dcache_tlb_cmd_put_partial  ? ~ dcache_tlb_ppp_array_if_cached :7'h0)|( dcache_tlb_cmd_amo_logical  ? ~ dcache_tlb_pal_array_if_cached :7'h0)|( dcache_tlb_cmd_amo_arithmetic  ? ~ dcache_tlb_paa_array_if_cached :7'h0); 
    wire[6:0] dcache_tlb_must_alloc_array =( dcache_tlb_cmd_put_partial  ? ~ dcache_tlb_ppp_array :7'h0)|( dcache_tlb_cmd_amo_logical  ? ~ dcache_tlb_pal_array :7'h0)|( dcache_tlb_cmd_amo_arithmetic  ? ~ dcache_tlb_paa_array :7'h0)|{7{ dcache_tlb_cmd_lrsc }}; 
    wire[6:0] dcache_tlb_pf_ld_array = dcache_tlb_cmd_read  ? (~ dcache_tlb_r_array &~ dcache_tlb_ptw_ae_array | dcache_tlb_ptw_pf_array )&~ dcache_tlb_ptw_gf_array :7'h0; 
    wire[6:0] dcache_tlb_pf_st_array = dcache_tlb_cmd_write_perms  ? (~ dcache_tlb_w_array &~ dcache_tlb_ptw_ae_array | dcache_tlb_ptw_pf_array )&~ dcache_tlb_ptw_gf_array :7'h0; 
    wire[6:0] dcache_tlb_pf_inst_array =(~ dcache_tlb_x_array &~ dcache_tlb_ptw_ae_array | dcache_tlb_ptw_pf_array )&~ dcache_tlb_ptw_gf_array ; 
    wire[1:0] dcache_tlb_lo ={ dcache_tlb_superpage_hits_1 , dcache_tlb_superpage_hits_0 }; 
    wire[1:0] dcache_tlb_lo_1 = dcache_tlb_lo ; 
    wire[1:0] dcache_tlb_hi ={ dcache_tlb_superpage_hits_3 , dcache_tlb_superpage_hits_2 }; 
    wire[1:0] dcache_tlb_hi_1 = dcache_tlb_hi ; 
    wire[1:0] dcache_tlb_state_reg_touch_way_sized ={| dcache_tlb_hi_1 , dcache_tlb_hi_1 [1]| dcache_tlb_lo_1 [1]}; 
    wire dcache_tlb_state_reg_set_left_older =~( dcache_tlb_state_reg_touch_way_sized [1]); 
    wire[1:0] dcache_tlb_state_reg_hi ={ dcache_tlb_state_reg_set_left_older ,~ dcache_tlb_state_reg_set_left_older &~( dcache_tlb_state_reg_touch_way_sized [0])}; 
    wire[20:0] dcache_tlb_io_resp_gpa_page ={1'h0, dcache_tlb_vpn }; 
    wire[19:0] dcache_pma_checker_vpn = dcache_s1_req_addr [31:12]; 
    wire[19:0] dcache_pma_checker_ppn = dcache_pma_checker_vpn ; 
    wire dcache_pma_checker_priv_s = dcache_s1_req_dprv [0]; 
    wire dcache_pma_checker_priv_uses_vm =~( dcache_s1_req_dprv [1]); 
    wire[19:0] dcache_pma_checker_mpu_ppn = dcache_s1_req_addr [31:12]; 
    wire[11:0] dcache_pma_checker_io_resp_gpa_offset = dcache_s1_req_addr [11:0]; 
    wire[31:0] dcache_pma_checker_mpu_physaddr ={ dcache_pma_checker_mpu_ppn , dcache_pma_checker_io_resp_gpa_offset }; 
    wire[2:0] dcache_pma_checker_mpu_priv ={1'h0, dcache_s1_req_dprv }; 
    wire[19:0] dcache__GEN_25 ={ dcache_pma_checker_mpu_physaddr [31:14],~( dcache_pma_checker_mpu_physaddr [13:12])}; 
    wire[5:0] dcache__GEN_26 ={ dcache_pma_checker_mpu_physaddr [31:28],~( dcache_pma_checker_mpu_physaddr [27:26])}; 
    wire[9:0] dcache__GEN_27 = dcache_pma_checker_mpu_physaddr [25:16]^10'h200; 
    wire[15:0] dcache__GEN_28 ={ dcache_pma_checker_mpu_physaddr [31:26], dcache__GEN_27 }; 
    wire dcache__GEN_29 = dcache_pma_checker_mpu_physaddr [31:14]!=18'h20000; 
    wire[15:0] dcache__GEN_30 ={ dcache_pma_checker_mpu_physaddr [31:17],~( dcache_pma_checker_mpu_physaddr [16])}; 
    wire[2:0] dcache__GEN_31 ={ dcache_pma_checker_mpu_physaddr [31],~( dcache_pma_checker_mpu_physaddr [30:29])}; 
    wire dcache_pma_checker_legal_address =~(| dcache__GEN_25 )|~(| dcache__GEN_26 )|~(| dcache__GEN_28 )|~ dcache__GEN_29 |~(|( dcache_pma_checker_mpu_physaddr [31:12]))|~(| dcache__GEN_30 )|~(| dcache__GEN_31 ); 
    wire dcache_pma_checker_homogeneous =~(|( dcache_pma_checker_mpu_physaddr [31:12]))|~(| dcache__GEN_25 )|~(| dcache__GEN_30 )|~(| dcache__GEN_28 )|~(| dcache__GEN_26 )|~(| dcache__GEN_31 )|~ dcache__GEN_29 ; 
    wire dcache_pma_checker_deny_access_to_debug =~( dcache_pma_checker_mpu_priv [2])&~(|( dcache_pma_checker_mpu_physaddr [31:12])); 
    wire dcache_pma_checker_prot_r = dcache_pma_checker_legal_address &~ dcache_pma_checker_deny_access_to_debug & dcache__pma_checker_pmp_io_r ; 
    wire dcache_pma_checker_newEntry_pr = dcache_pma_checker_prot_r ; 
    wire[2:0] dcache__GEN_32 ={ dcache_pma_checker_mpu_physaddr [30], dcache_pma_checker_mpu_physaddr [27], dcache_pma_checker_mpu_physaddr [16]}; 
    wire[2:0] dcache__GEN_33 ={ dcache_pma_checker_mpu_physaddr [31:30],~( dcache_pma_checker_mpu_physaddr [27])}; 
    wire[1:0] dcache__GEN_34 ={ dcache_pma_checker_mpu_physaddr [31],~( dcache_pma_checker_mpu_physaddr [30])}; 
    wire dcache_pma_checker_prot_w = dcache_pma_checker_legal_address &(~(| dcache__GEN_32 )|~(| dcache__GEN_33 )|~(| dcache__GEN_34 ))&~ dcache_pma_checker_deny_access_to_debug & dcache__pma_checker_pmp_io_w ; 
    wire dcache_pma_checker_newEntry_pw = dcache_pma_checker_prot_w ; 
    wire dcache_pma_checker_prot_pp = dcache_pma_checker_legal_address &(~(| dcache__GEN_32 )|~(| dcache__GEN_33 )|~(| dcache__GEN_34 )); 
    wire dcache_pma_checker_newEntry_ppp = dcache_pma_checker_prot_pp ; 
    wire dcache_pma_checker_prot_al = dcache_pma_checker_legal_address &(~(| dcache__GEN_32 )|~(| dcache__GEN_33 )); 
    wire dcache_pma_checker_newEntry_pal = dcache_pma_checker_prot_al ; 
    wire dcache_pma_checker_prot_aa = dcache_pma_checker_legal_address &(~(| dcache__GEN_32 )|~(| dcache__GEN_33 )); 
    wire dcache_pma_checker_newEntry_paa = dcache_pma_checker_prot_aa ; 
    wire dcache_pma_checker_prot_x = dcache_pma_checker_legal_address &({ dcache_pma_checker_mpu_physaddr [30], dcache_pma_checker_mpu_physaddr [27], dcache_pma_checker_mpu_physaddr [25]}==3'h0|~(| dcache__GEN_34 ))&~ dcache_pma_checker_deny_access_to_debug & dcache__pma_checker_pmp_io_x ; 
    wire dcache_pma_checker_newEntry_px = dcache_pma_checker_prot_x ; 
    wire dcache_pma_checker_prot_eff = dcache_pma_checker_legal_address &({ dcache_pma_checker_mpu_physaddr [31:30], dcache_pma_checker_mpu_physaddr [27], dcache_pma_checker_mpu_physaddr [25], dcache_pma_checker_mpu_physaddr [16], dcache_pma_checker_mpu_physaddr [13]}==6'h0|{ dcache_pma_checker_mpu_physaddr [31:30], dcache_pma_checker_mpu_physaddr [27], dcache__GEN_27 [9], dcache_pma_checker_mpu_physaddr [16]}==5'h0|~(| dcache__GEN_33 )|~(| dcache__GEN_34 )); 
    wire dcache_pma_checker_newEntry_eff = dcache_pma_checker_prot_eff ; 
    wire[1:0] dcache_pma_checker_hitsVec_idx = dcache_pma_checker_vpn [1:0]; 
    wire[1:0] dcache__GEN_35 ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_lo_hi_hi ; 
  assign  dcache_pma_checker_special_entry_data_0_lo_lo_hi_hi = dcache__GEN_35 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi_hi = dcache__GEN_35 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi_hi = dcache__GEN_35 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi_hi = dcache__GEN_35 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi_hi = dcache__GEN_35 ; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi_hi ; 
  assign  dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi_hi = dcache__GEN_35 ; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_lo_lo_hi ={ dcache_pma_checker_special_entry_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_special_entry_data_0_lo_lo ={ dcache_pma_checker_special_entry_data_0_lo_lo_hi ,2'h0}; 
    wire[1:0] dcache__GEN_36 ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_hi_lo_hi ; 
  assign  dcache_pma_checker_special_entry_data_0_lo_hi_lo_hi = dcache__GEN_36 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo_hi ; 
  assign  dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo_hi = dcache__GEN_36 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo_hi ; 
  assign  dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo_hi = dcache__GEN_36 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo_hi ; 
  assign  dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo_hi = dcache__GEN_36 ; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo_hi ; 
  assign  dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo_hi = dcache__GEN_36 ; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo_hi ; 
  assign  dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo_hi = dcache__GEN_36 ; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_lo_hi_lo ={ dcache_pma_checker_special_entry_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[2:0] dcache__GEN_37 ={2'h0, dcache_pma_checker_newEntry_pw }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_lo_hi_hi ; 
  assign  dcache_pma_checker_special_entry_data_0_lo_hi_hi = dcache__GEN_37 ; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi = dcache__GEN_37 ; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi = dcache__GEN_37 ; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi = dcache__GEN_37 ; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi ; 
  assign  dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi = dcache__GEN_37 ; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi ; 
  assign  dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi = dcache__GEN_37 ; 
    wire[5:0] dcache_pma_checker_special_entry_data_0_lo_hi ={ dcache_pma_checker_special_entry_data_0_lo_hi_hi , dcache_pma_checker_special_entry_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_special_entry_data_0_lo ={ dcache_pma_checker_special_entry_data_0_lo_hi , dcache_pma_checker_special_entry_data_0_lo_lo }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[5:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_0_data_0_lo ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi , dcache_pma_checker_superpage_entries_0_data_0_lo_lo }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[5:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_1_data_0_lo ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi , dcache_pma_checker_superpage_entries_1_data_0_lo_lo }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[5:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_2_data_0_lo ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi , dcache_pma_checker_superpage_entries_2_data_0_lo_lo }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[5:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_3_data_0_lo ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi , dcache_pma_checker_superpage_entries_3_data_0_lo_lo }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi ={ dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo ={ dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi ,2'h0}; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[5:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi , dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_sectored_entries_0_0_data_lo ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi , dcache_pma_checker_sectored_entries_0_0_data_lo_lo }; 
    wire[1:0] dcache_pma_checker_ptw_ae_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_ae_ptw , dcache__pma_checker_entries_barrier_1_io_y_ae_ptw }; 
    wire[2:0] dcache_pma_checker_ptw_ae_array_lo ={ dcache_pma_checker_ptw_ae_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_ae_ptw }; 
    wire[1:0] dcache_pma_checker_ptw_ae_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_ae_ptw , dcache__pma_checker_entries_barrier_4_io_y_ae_ptw }; 
    wire[2:0] dcache_pma_checker_ptw_ae_array_hi ={ dcache_pma_checker_ptw_ae_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_ae_ptw }; 
    wire[6:0] dcache_pma_checker_ptw_ae_array ={1'h0, dcache_pma_checker_ptw_ae_array_hi , dcache_pma_checker_ptw_ae_array_lo }; 
    wire[1:0] dcache_pma_checker_final_ae_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_ae_final , dcache__pma_checker_entries_barrier_1_io_y_ae_final }; 
    wire[2:0] dcache_pma_checker_final_ae_array_lo ={ dcache_pma_checker_final_ae_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_ae_final }; 
    wire[1:0] dcache_pma_checker_final_ae_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_ae_final , dcache__pma_checker_entries_barrier_4_io_y_ae_final }; 
    wire[2:0] dcache_pma_checker_final_ae_array_hi ={ dcache_pma_checker_final_ae_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_ae_final }; 
    wire[6:0] dcache_pma_checker_final_ae_array ={1'h0, dcache_pma_checker_final_ae_array_hi , dcache_pma_checker_final_ae_array_lo }; 
    wire[1:0] dcache_pma_checker_ptw_pf_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_pf , dcache__pma_checker_entries_barrier_1_io_y_pf }; 
    wire[2:0] dcache_pma_checker_ptw_pf_array_lo ={ dcache_pma_checker_ptw_pf_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_pf }; 
    wire[1:0] dcache_pma_checker_ptw_pf_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_pf , dcache__pma_checker_entries_barrier_4_io_y_pf }; 
    wire[2:0] dcache_pma_checker_ptw_pf_array_hi ={ dcache_pma_checker_ptw_pf_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_pf }; 
    wire[6:0] dcache_pma_checker_ptw_pf_array ={1'h0, dcache_pma_checker_ptw_pf_array_hi , dcache_pma_checker_ptw_pf_array_lo }; 
    wire[1:0] dcache_pma_checker_ptw_gf_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_gf , dcache__pma_checker_entries_barrier_1_io_y_gf }; 
    wire[2:0] dcache_pma_checker_ptw_gf_array_lo ={ dcache_pma_checker_ptw_gf_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_gf }; 
    wire[1:0] dcache_pma_checker_ptw_gf_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_gf , dcache__pma_checker_entries_barrier_4_io_y_gf }; 
    wire[2:0] dcache_pma_checker_ptw_gf_array_hi ={ dcache_pma_checker_ptw_gf_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_gf }; 
    wire[6:0] dcache_pma_checker_ptw_gf_array ={1'h0, dcache_pma_checker_ptw_gf_array_hi , dcache_pma_checker_ptw_gf_array_lo }; 
    wire[1:0] dcache__GEN_38 ={ dcache__pma_checker_entries_barrier_2_io_y_u , dcache__pma_checker_entries_barrier_1_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_lo_hi ; 
  assign  dcache_pma_checker_priv_rw_ok_lo_hi = dcache__GEN_38 ; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_lo_hi_1 ; 
  assign  dcache_pma_checker_priv_rw_ok_lo_hi_1 = dcache__GEN_38 ; 
    wire[1:0] dcache_pma_checker_priv_x_ok_lo_hi ; 
  assign  dcache_pma_checker_priv_x_ok_lo_hi = dcache__GEN_38 ; 
    wire[1:0] dcache_pma_checker_priv_x_ok_lo_hi_1 ; 
  assign  dcache_pma_checker_priv_x_ok_lo_hi_1 = dcache__GEN_38 ; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_lo ={ dcache_pma_checker_priv_rw_ok_lo_hi , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[1:0] dcache__GEN_39 ={ dcache__pma_checker_entries_barrier_5_io_y_u , dcache__pma_checker_entries_barrier_4_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_hi_hi ; 
  assign  dcache_pma_checker_priv_rw_ok_hi_hi = dcache__GEN_39 ; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_hi_hi_1 ; 
  assign  dcache_pma_checker_priv_rw_ok_hi_hi_1 = dcache__GEN_39 ; 
    wire[1:0] dcache_pma_checker_priv_x_ok_hi_hi ; 
  assign  dcache_pma_checker_priv_x_ok_hi_hi = dcache__GEN_39 ; 
    wire[1:0] dcache_pma_checker_priv_x_ok_hi_hi_1 ; 
  assign  dcache_pma_checker_priv_x_ok_hi_hi_1 = dcache__GEN_39 ; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_hi ={ dcache_pma_checker_priv_rw_ok_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_lo_1 ={ dcache_pma_checker_priv_rw_ok_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_hi_1 ={ dcache_pma_checker_priv_rw_ok_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_pma_checker_priv_rw_ok =( dcache_pma_checker_priv_s  ? 6'h0:{ dcache_pma_checker_priv_rw_ok_hi , dcache_pma_checker_priv_rw_ok_lo })|( dcache_pma_checker_priv_s  ? ~{ dcache_pma_checker_priv_rw_ok_hi_1 , dcache_pma_checker_priv_rw_ok_lo_1 }:6'h0); 
    wire[2:0] dcache_pma_checker_priv_x_ok_lo ={ dcache_pma_checker_priv_x_ok_lo_hi , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_hi ={ dcache_pma_checker_priv_x_ok_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_lo_1 ={ dcache_pma_checker_priv_x_ok_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_hi_1 ={ dcache_pma_checker_priv_x_ok_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_pma_checker_priv_x_ok = dcache_pma_checker_priv_s  ? ~{ dcache_pma_checker_priv_x_ok_hi , dcache_pma_checker_priv_x_ok_lo }:{ dcache_pma_checker_priv_x_ok_hi_1 , dcache_pma_checker_priv_x_ok_lo_1 }; 
    wire[1:0] dcache_pma_checker_stage1_bypass_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_ae_stage2 , dcache__pma_checker_entries_barrier_1_io_y_ae_stage2 }; 
    wire[2:0] dcache_pma_checker_stage1_bypass_lo ={ dcache_pma_checker_stage1_bypass_lo_hi , dcache__pma_checker_entries_barrier_io_y_ae_stage2 }; 
    wire[1:0] dcache_pma_checker_stage1_bypass_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_ae_stage2 , dcache__pma_checker_entries_barrier_4_io_y_ae_stage2 }; 
    wire[2:0] dcache_pma_checker_stage1_bypass_hi ={ dcache_pma_checker_stage1_bypass_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_ae_stage2 }; 
    wire[1:0] dcache_pma_checker_r_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_sr , dcache__pma_checker_entries_barrier_1_io_y_sr }; 
    wire[2:0] dcache_pma_checker_r_array_lo ={ dcache_pma_checker_r_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_sr }; 
    wire[1:0] dcache_pma_checker_r_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_sr , dcache__pma_checker_entries_barrier_4_io_y_sr }; 
    wire[2:0] dcache_pma_checker_r_array_hi ={ dcache_pma_checker_r_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_sr }; 
    wire[1:0] dcache__GEN_40 ={ dcache__pma_checker_entries_barrier_2_io_y_sx , dcache__pma_checker_entries_barrier_1_io_y_sx }; 
    wire[1:0] dcache_pma_checker_r_array_lo_hi_1 ; 
  assign  dcache_pma_checker_r_array_lo_hi_1 = dcache__GEN_40 ; 
    wire[1:0] dcache_pma_checker_x_array_lo_hi ; 
  assign  dcache_pma_checker_x_array_lo_hi = dcache__GEN_40 ; 
    wire[2:0] dcache_pma_checker_r_array_lo_1 ={ dcache_pma_checker_r_array_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_sx }; 
    wire[1:0] dcache__GEN_41 ={ dcache__pma_checker_entries_barrier_5_io_y_sx , dcache__pma_checker_entries_barrier_4_io_y_sx }; 
    wire[1:0] dcache_pma_checker_r_array_hi_hi_1 ; 
  assign  dcache_pma_checker_r_array_hi_hi_1 = dcache__GEN_41 ; 
    wire[1:0] dcache_pma_checker_x_array_hi_hi ; 
  assign  dcache_pma_checker_x_array_hi_hi = dcache__GEN_41 ; 
    wire[2:0] dcache_pma_checker_r_array_hi_1 ={ dcache_pma_checker_r_array_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_pma_checker_r_array ={1'h1, dcache_pma_checker_priv_rw_ok &{ dcache_pma_checker_r_array_hi , dcache_pma_checker_r_array_lo }}; 
    wire[1:0] dcache_pma_checker_w_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_sw , dcache__pma_checker_entries_barrier_1_io_y_sw }; 
    wire[2:0] dcache_pma_checker_w_array_lo ={ dcache_pma_checker_w_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_sw }; 
    wire[1:0] dcache_pma_checker_w_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_sw , dcache__pma_checker_entries_barrier_4_io_y_sw }; 
    wire[2:0] dcache_pma_checker_w_array_hi ={ dcache_pma_checker_w_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_sw }; 
    wire[6:0] dcache_pma_checker_w_array ={1'h1, dcache_pma_checker_priv_rw_ok &{ dcache_pma_checker_w_array_hi , dcache_pma_checker_w_array_lo }}; 
    wire[2:0] dcache_pma_checker_x_array_lo ={ dcache_pma_checker_x_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_sx }; 
    wire[2:0] dcache_pma_checker_x_array_hi ={ dcache_pma_checker_x_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_pma_checker_x_array ={1'h1, dcache_pma_checker_priv_x_ok &{ dcache_pma_checker_x_array_hi , dcache_pma_checker_x_array_lo }}; 
    wire[1:0] dcache_pma_checker_hr_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_hr , dcache__pma_checker_entries_barrier_1_io_y_hr }; 
    wire[2:0] dcache_pma_checker_hr_array_lo ={ dcache_pma_checker_hr_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_hr }; 
    wire[1:0] dcache_pma_checker_hr_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_hr , dcache__pma_checker_entries_barrier_4_io_y_hr }; 
    wire[2:0] dcache_pma_checker_hr_array_hi ={ dcache_pma_checker_hr_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_hr }; 
    wire[1:0] dcache__GEN_42 ={ dcache__pma_checker_entries_barrier_2_io_y_hx , dcache__pma_checker_entries_barrier_1_io_y_hx }; 
    wire[1:0] dcache_pma_checker_hr_array_lo_hi_1 ; 
  assign  dcache_pma_checker_hr_array_lo_hi_1 = dcache__GEN_42 ; 
    wire[1:0] dcache_pma_checker_hx_array_lo_hi ; 
  assign  dcache_pma_checker_hx_array_lo_hi = dcache__GEN_42 ; 
    wire[2:0] dcache_pma_checker_hr_array_lo_1 ={ dcache_pma_checker_hr_array_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_hx }; 
    wire[1:0] dcache__GEN_43 ={ dcache__pma_checker_entries_barrier_5_io_y_hx , dcache__pma_checker_entries_barrier_4_io_y_hx }; 
    wire[1:0] dcache_pma_checker_hr_array_hi_hi_1 ; 
  assign  dcache_pma_checker_hr_array_hi_hi_1 = dcache__GEN_43 ; 
    wire[1:0] dcache_pma_checker_hx_array_hi_hi ; 
  assign  dcache_pma_checker_hx_array_hi_hi = dcache__GEN_43 ; 
    wire[2:0] dcache_pma_checker_hr_array_hi_1 ={ dcache_pma_checker_hr_array_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_hx }; 
    wire[1:0] dcache_pma_checker_hw_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_hw , dcache__pma_checker_entries_barrier_1_io_y_hw }; 
    wire[2:0] dcache_pma_checker_hw_array_lo ={ dcache_pma_checker_hw_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_hw }; 
    wire[1:0] dcache_pma_checker_hw_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_hw , dcache__pma_checker_entries_barrier_4_io_y_hw }; 
    wire[2:0] dcache_pma_checker_hw_array_hi ={ dcache_pma_checker_hw_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_hw }; 
    wire[2:0] dcache_pma_checker_hx_array_lo ={ dcache_pma_checker_hx_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_hx }; 
    wire[2:0] dcache_pma_checker_hx_array_hi ={ dcache_pma_checker_hx_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_hx }; 
    wire[1:0] dcache_pma_checker_pr_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_pr , dcache__pma_checker_entries_barrier_io_y_pr }; 
    wire[1:0] dcache_pma_checker_pr_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_pr , dcache__pma_checker_entries_barrier_3_io_y_pr }; 
    wire[2:0] dcache_pma_checker_pr_array_hi ={ dcache_pma_checker_pr_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_pr }; 
    wire[6:0] dcache_pma_checker__pr_array_T_4 = dcache_pma_checker_ptw_ae_array | dcache_pma_checker_final_ae_array ; 
    wire[6:0] dcache_pma_checker_pr_array ={{2{ dcache_pma_checker_prot_r }}, dcache_pma_checker_pr_array_hi , dcache_pma_checker_pr_array_lo }&~ dcache_pma_checker__pr_array_T_4 ; 
    wire[1:0] dcache_pma_checker_pw_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_pw , dcache__pma_checker_entries_barrier_io_y_pw }; 
    wire[1:0] dcache_pma_checker_pw_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_pw , dcache__pma_checker_entries_barrier_3_io_y_pw }; 
    wire[2:0] dcache_pma_checker_pw_array_hi ={ dcache_pma_checker_pw_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_pw }; 
    wire[6:0] dcache_pma_checker_pw_array ={{2{ dcache_pma_checker_prot_w }}, dcache_pma_checker_pw_array_hi , dcache_pma_checker_pw_array_lo }&~ dcache_pma_checker__pr_array_T_4 ; 
    wire[1:0] dcache_pma_checker_px_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_px , dcache__pma_checker_entries_barrier_io_y_px }; 
    wire[1:0] dcache_pma_checker_px_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_px , dcache__pma_checker_entries_barrier_3_io_y_px }; 
    wire[2:0] dcache_pma_checker_px_array_hi ={ dcache_pma_checker_px_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_px }; 
    wire[6:0] dcache_pma_checker_px_array ={{2{ dcache_pma_checker_prot_x }}, dcache_pma_checker_px_array_hi , dcache_pma_checker_px_array_lo }&~ dcache_pma_checker__pr_array_T_4 ; 
    wire[1:0] dcache_pma_checker_eff_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_eff , dcache__pma_checker_entries_barrier_io_y_eff }; 
    wire[1:0] dcache_pma_checker_eff_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_eff , dcache__pma_checker_entries_barrier_3_io_y_eff }; 
    wire[2:0] dcache_pma_checker_eff_array_hi ={ dcache_pma_checker_eff_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_eff }; 
    wire[6:0] dcache_pma_checker_eff_array ={{2{ dcache_pma_checker_prot_eff }}, dcache_pma_checker_eff_array_hi , dcache_pma_checker_eff_array_lo }; 
    wire[1:0] dcache__GEN_44 ={ dcache__pma_checker_entries_barrier_1_io_y_c , dcache__pma_checker_entries_barrier_io_y_c }; 
    wire[1:0] dcache_pma_checker_c_array_lo ; 
  assign  dcache_pma_checker_c_array_lo = dcache__GEN_44 ; 
    wire[1:0] dcache_pma_checker_prefetchable_array_lo ; 
  assign  dcache_pma_checker_prefetchable_array_lo = dcache__GEN_44 ; 
    wire[1:0] dcache__GEN_45 ={ dcache__pma_checker_entries_barrier_4_io_y_c , dcache__pma_checker_entries_barrier_3_io_y_c }; 
    wire[1:0] dcache_pma_checker_c_array_hi_hi ; 
  assign  dcache_pma_checker_c_array_hi_hi = dcache__GEN_45 ; 
    wire[1:0] dcache_pma_checker_prefetchable_array_hi_hi ; 
  assign  dcache_pma_checker_prefetchable_array_hi_hi = dcache__GEN_45 ; 
    wire[2:0] dcache_pma_checker_c_array_hi ={ dcache_pma_checker_c_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_pma_checker_c_array ={2'h0, dcache_pma_checker_c_array_hi , dcache_pma_checker_c_array_lo }; 
    wire[1:0] dcache_pma_checker_ppp_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_ppp , dcache__pma_checker_entries_barrier_io_y_ppp }; 
    wire[1:0] dcache_pma_checker_ppp_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_ppp , dcache__pma_checker_entries_barrier_3_io_y_ppp }; 
    wire[2:0] dcache_pma_checker_ppp_array_hi ={ dcache_pma_checker_ppp_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_ppp }; 
    wire[6:0] dcache_pma_checker_ppp_array ={{2{ dcache_pma_checker_prot_pp }}, dcache_pma_checker_ppp_array_hi , dcache_pma_checker_ppp_array_lo }; 
    wire[1:0] dcache_pma_checker_paa_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_paa , dcache__pma_checker_entries_barrier_io_y_paa }; 
    wire[1:0] dcache_pma_checker_paa_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_paa , dcache__pma_checker_entries_barrier_3_io_y_paa }; 
    wire[2:0] dcache_pma_checker_paa_array_hi ={ dcache_pma_checker_paa_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_paa }; 
    wire[6:0] dcache_pma_checker_paa_array ={{2{ dcache_pma_checker_prot_aa }}, dcache_pma_checker_paa_array_hi , dcache_pma_checker_paa_array_lo }; 
    wire[1:0] dcache_pma_checker_pal_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_pal , dcache__pma_checker_entries_barrier_io_y_pal }; 
    wire[1:0] dcache_pma_checker_pal_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_pal , dcache__pma_checker_entries_barrier_3_io_y_pal }; 
    wire[2:0] dcache_pma_checker_pal_array_hi ={ dcache_pma_checker_pal_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_pal }; 
    wire[6:0] dcache_pma_checker_pal_array ={{2{ dcache_pma_checker_prot_al }}, dcache_pma_checker_pal_array_hi , dcache_pma_checker_pal_array_lo }; 
    wire[6:0] dcache_pma_checker_ppp_array_if_cached = dcache_pma_checker_ppp_array | dcache_pma_checker_c_array ; 
    wire[6:0] dcache_pma_checker_paa_array_if_cached = dcache_pma_checker_paa_array | dcache_pma_checker_c_array ; 
    wire[6:0] dcache_pma_checker_pal_array_if_cached = dcache_pma_checker_pal_array | dcache_pma_checker_c_array ; 
    wire[2:0] dcache_pma_checker_prefetchable_array_hi ={ dcache_pma_checker_prefetchable_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_pma_checker_prefetchable_array ={2'h0, dcache_pma_checker_prefetchable_array_hi , dcache_pma_checker_prefetchable_array_lo }; 
    wire dcache_pma_checker_misaligned =|( dcache_s1_req_addr [3:0]&(4'h1<< dcache_s1_req_size )-4'h1); 
    wire dcache_pma_checker__cmd_lrsc_T = dcache_s1_req_cmd ==5'h6; 
    wire dcache_pma_checker__cmd_lrsc_T_1 = dcache_s1_req_cmd ==5'h7; 
    wire dcache_pma_checker_cmd_lrsc = dcache_pma_checker__cmd_lrsc_T | dcache_pma_checker__cmd_lrsc_T_1 ; 
    wire dcache_pma_checker__cmd_read_T_7 = dcache_s1_req_cmd ==5'h4; 
    wire dcache_pma_checker__cmd_read_T_8 = dcache_s1_req_cmd ==5'h9; 
    wire dcache_pma_checker__cmd_read_T_9 = dcache_s1_req_cmd ==5'hA; 
    wire dcache_pma_checker__cmd_read_T_10 = dcache_s1_req_cmd ==5'hB; 
    wire dcache_pma_checker_cmd_amo_logical = dcache_pma_checker__cmd_read_T_7 | dcache_pma_checker__cmd_read_T_8 | dcache_pma_checker__cmd_read_T_9 | dcache_pma_checker__cmd_read_T_10 ; 
    wire dcache_pma_checker__cmd_read_T_14 = dcache_s1_req_cmd ==5'h8; 
    wire dcache_pma_checker__cmd_read_T_15 = dcache_s1_req_cmd ==5'hC; 
    wire dcache_pma_checker__cmd_read_T_16 = dcache_s1_req_cmd ==5'hD; 
    wire dcache_pma_checker__cmd_read_T_17 = dcache_s1_req_cmd ==5'hE; 
    wire dcache_pma_checker__cmd_read_T_18 = dcache_s1_req_cmd ==5'hF; 
    wire dcache_pma_checker_cmd_amo_arithmetic = dcache_pma_checker__cmd_read_T_14 | dcache_pma_checker__cmd_read_T_15 | dcache_pma_checker__cmd_read_T_16 | dcache_pma_checker__cmd_read_T_17 | dcache_pma_checker__cmd_read_T_18 ; 
    wire dcache_pma_checker_cmd_put_partial = dcache_s1_req_cmd ==5'h11; 
    wire dcache_pma_checker_cmd_read = dcache_s1_req_cmd ==5'h0| dcache_s1_req_cmd ==5'h10| dcache_pma_checker__cmd_lrsc_T | dcache_pma_checker__cmd_lrsc_T_1 | dcache_pma_checker__cmd_read_T_7 | dcache_pma_checker__cmd_read_T_8 | dcache_pma_checker__cmd_read_T_9 | dcache_pma_checker__cmd_read_T_10 | dcache_pma_checker__cmd_read_T_14 | dcache_pma_checker__cmd_read_T_15 | dcache_pma_checker__cmd_read_T_16 | dcache_pma_checker__cmd_read_T_17 | dcache_pma_checker__cmd_read_T_18 ; 
    wire dcache_pma_checker_cmd_write = dcache_s1_req_cmd ==5'h1| dcache_pma_checker_cmd_put_partial | dcache_pma_checker__cmd_lrsc_T_1 | dcache_pma_checker__cmd_read_T_7 | dcache_pma_checker__cmd_read_T_8 | dcache_pma_checker__cmd_read_T_9 | dcache_pma_checker__cmd_read_T_10 | dcache_pma_checker__cmd_read_T_14 | dcache_pma_checker__cmd_read_T_15 | dcache_pma_checker__cmd_read_T_16 | dcache_pma_checker__cmd_read_T_17 | dcache_pma_checker__cmd_read_T_18 ; 
    wire dcache_pma_checker_cmd_write_perms = dcache_pma_checker_cmd_write | dcache_s1_req_cmd ==5'h5| dcache_s1_req_cmd ==5'h17; 
    wire[6:0] dcache_pma_checker_ae_array =( dcache_pma_checker_misaligned  ?  dcache_pma_checker_eff_array :7'h0)|{7{ dcache_pma_checker_cmd_lrsc }}; 
    wire[6:0] dcache_pma_checker_ae_ld_array = dcache_pma_checker_cmd_read  ?  dcache_pma_checker_ae_array |~ dcache_pma_checker_pr_array :7'h0; 
    wire[6:0] dcache_pma_checker_ae_st_array =( dcache_pma_checker_cmd_write_perms  ?  dcache_pma_checker_ae_array |~ dcache_pma_checker_pw_array :7'h0)|( dcache_pma_checker_cmd_put_partial  ? ~ dcache_pma_checker_ppp_array_if_cached :7'h0)|( dcache_pma_checker_cmd_amo_logical  ? ~ dcache_pma_checker_pal_array_if_cached :7'h0)|( dcache_pma_checker_cmd_amo_arithmetic  ? ~ dcache_pma_checker_paa_array_if_cached :7'h0); 
    wire[6:0] dcache_pma_checker_must_alloc_array =( dcache_pma_checker_cmd_put_partial  ? ~ dcache_pma_checker_ppp_array :7'h0)|( dcache_pma_checker_cmd_amo_logical  ? ~ dcache_pma_checker_pal_array :7'h0)|( dcache_pma_checker_cmd_amo_arithmetic  ? ~ dcache_pma_checker_paa_array :7'h0)|{7{ dcache_pma_checker_cmd_lrsc }}; 
    wire[6:0] dcache_pma_checker_pf_ld_array = dcache_pma_checker_cmd_read  ? (~ dcache_pma_checker_r_array &~ dcache_pma_checker_ptw_ae_array | dcache_pma_checker_ptw_pf_array )&~ dcache_pma_checker_ptw_gf_array :7'h0; 
    wire[6:0] dcache_pma_checker_pf_st_array = dcache_pma_checker_cmd_write_perms  ? (~ dcache_pma_checker_w_array &~ dcache_pma_checker_ptw_ae_array | dcache_pma_checker_ptw_pf_array )&~ dcache_pma_checker_ptw_gf_array :7'h0; 
    wire[6:0] dcache_pma_checker_pf_inst_array =(~ dcache_pma_checker_x_array &~ dcache_pma_checker_ptw_ae_array | dcache_pma_checker_ptw_pf_array )&~ dcache_pma_checker_ptw_gf_array ; 
    wire[1:0] dcache_pma_checker_lo ={ dcache_pma_checker_superpage_hits_1 , dcache_pma_checker_superpage_hits_0 }; 
    wire[1:0] dcache_pma_checker_lo_1 = dcache_pma_checker_lo ; 
    wire[1:0] dcache_pma_checker_hi ={ dcache_pma_checker_superpage_hits_3 , dcache_pma_checker_superpage_hits_2 }; 
    wire[1:0] dcache_pma_checker_hi_1 = dcache_pma_checker_hi ; 
    wire[1:0] dcache_pma_checker_state_reg_touch_way_sized ={| dcache_pma_checker_hi_1 , dcache_pma_checker_hi_1 [1]| dcache_pma_checker_lo_1 [1]}; 
    wire dcache_pma_checker_state_reg_set_left_older =~( dcache_pma_checker_state_reg_touch_way_sized [1]); 
    wire[1:0] dcache_pma_checker_state_reg_hi ={ dcache_pma_checker_state_reg_set_left_older ,~ dcache_pma_checker_state_reg_set_left_older &~( dcache_pma_checker_state_reg_touch_way_sized [0])}; 
    wire[20:0] dcache_pma_checker_io_resp_gpa_page ={1'h0, dcache_pma_checker_vpn }; 
    wire[1:0] dcache_lfsr_lo_lo_lo ={ dcache__lfsr_prng_io_out_1 , dcache__lfsr_prng_io_out_0 }; 
    wire[1:0] dcache_lfsr_lo_lo_hi ={ dcache__lfsr_prng_io_out_3 , dcache__lfsr_prng_io_out_2 }; 
    wire[3:0] dcache_lfsr_lo_lo ={ dcache_lfsr_lo_lo_hi , dcache_lfsr_lo_lo_lo }; 
    wire[1:0] dcache_lfsr_lo_hi_lo ={ dcache__lfsr_prng_io_out_5 , dcache__lfsr_prng_io_out_4 }; 
    wire[1:0] dcache_lfsr_lo_hi_hi ={ dcache__lfsr_prng_io_out_7 , dcache__lfsr_prng_io_out_6 }; 
    wire[3:0] dcache_lfsr_lo_hi ={ dcache_lfsr_lo_hi_hi , dcache_lfsr_lo_hi_lo }; 
    wire[7:0] dcache_lfsr_lo ={ dcache_lfsr_lo_hi , dcache_lfsr_lo_lo }; 
    wire[1:0] dcache_lfsr_hi_lo_lo ={ dcache__lfsr_prng_io_out_9 , dcache__lfsr_prng_io_out_8 }; 
    wire[1:0] dcache_lfsr_hi_lo_hi ={ dcache__lfsr_prng_io_out_11 , dcache__lfsr_prng_io_out_10 }; 
    wire[3:0] dcache_lfsr_hi_lo ={ dcache_lfsr_hi_lo_hi , dcache_lfsr_hi_lo_lo }; 
    wire[1:0] dcache_lfsr_hi_hi_lo ={ dcache__lfsr_prng_io_out_13 , dcache__lfsr_prng_io_out_12 }; 
    wire[1:0] dcache_lfsr_hi_hi_hi ={ dcache__lfsr_prng_io_out_15 , dcache__lfsr_prng_io_out_14 }; 
    wire[3:0] dcache_lfsr_hi_hi ={ dcache_lfsr_hi_hi_hi , dcache_lfsr_hi_hi_lo }; 
    wire[7:0] dcache_lfsr_hi ={ dcache_lfsr_hi_hi , dcache_lfsr_hi_lo }; 
    wire[15:0] dcache_lfsr ={ dcache_lfsr_hi , dcache_lfsr_lo }; 
    wire[31:0] dcache_s2_vaddr ; 
    wire dcache_metaArb__grant_T_2 = dcache_metaArb_io_in_2_valid | dcache_metaArb_io_in_3_valid ; 
    wire dcache_metaArb_grant_3 =~ dcache_metaArb_io_in_2_valid ; 
    wire dcache_metaArb_grant_4 =~ dcache_metaArb__grant_T_2 ; 
    wire dcache_metaArb_grant_5 =~ dcache_metaArb__grant_T_2 ; 
    wire dcache_metaArb_grant_6 =~ dcache_metaArb__grant_T_2 ; 
    wire dcache_metaArb_grant_7 =~ dcache_metaArb__grant_T_2 ; 
    wire dcache__GEN_46 = dcache_dataArb_io_in_0_valid | dcache_dataArb_io_in_1_valid ; 
    wire dcache_pstore_drain ; 
    wire dcache_dataArb__grant_T = dcache_dataArb_io_in_0_valid | dcache_dataArb_io_in_1_valid ; 
    wire dcache_dataArb_grant_1 =~ dcache_dataArb_io_in_0_valid ; 
    wire dcache_dataArb_grant_2 =~ dcache_dataArb__grant_T ; 
    wire dcache_dataArb_grant_3 =~ dcache_dataArb__grant_T ; 
    wire dcache_dataArb_io_out_valid =~ dcache_dataArb_grant_3 | dcache_dataArb_io_in_3_valid ; 
  assign  dcache_nodeOut_a_deq_valid = dcache_tl_out_a_valid ; 
  assign  dcache_nodeOut_a_deq_bits_opcode = dcache_tl_out_a_bits_opcode ; 
  assign  dcache_nodeOut_a_deq_bits_param = dcache_tl_out_a_bits_param ; 
  assign  dcache_nodeOut_a_deq_bits_size = dcache_tl_out_a_bits_size ; 
  assign  dcache_nodeOut_a_deq_bits_address = dcache_tl_out_a_bits_address ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_bufferable = dcache_tl_out_a_bits_user_amba_prot_bufferable ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_modifiable = dcache_tl_out_a_bits_user_amba_prot_modifiable ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_readalloc = dcache_tl_out_a_bits_user_amba_prot_readalloc ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_writealloc = dcache_tl_out_a_bits_user_amba_prot_writealloc ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_privileged = dcache_tl_out_a_bits_user_amba_prot_privileged ; 
  assign  dcache_nodeOut_a_deq_bits_mask = dcache_tl_out_a_bits_mask ; 
  assign  dcache_nodeOut_a_deq_bits_data = dcache_tl_out_a_bits_data ; 
    wire dcache_tl_out_a_ready = dcache_nodeOut_a_deq_ready ; 
    wire dcache_nodeOut_a_valid = dcache_nodeOut_a_deq_valid ; 
    wire[2:0] dcache_nodeOut_a_bits_opcode = dcache_nodeOut_a_deq_bits_opcode ; 
    wire[2:0] dcache_nodeOut_a_bits_param = dcache_nodeOut_a_deq_bits_param ; 
    wire[3:0] dcache_nodeOut_a_bits_size = dcache_nodeOut_a_deq_bits_size ; 
    wire[31:0] dcache_nodeOut_a_bits_address = dcache_nodeOut_a_deq_bits_address ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_bufferable = dcache_nodeOut_a_deq_bits_user_amba_prot_bufferable ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_modifiable = dcache_nodeOut_a_deq_bits_user_amba_prot_modifiable ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_readalloc = dcache_nodeOut_a_deq_bits_user_amba_prot_readalloc ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_writealloc = dcache_nodeOut_a_deq_bits_user_amba_prot_writealloc ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_privileged = dcache_nodeOut_a_deq_bits_user_amba_prot_privileged ; 
    wire[3:0] dcache_nodeOut_a_bits_mask = dcache_nodeOut_a_deq_bits_mask ; 
    wire[31:0] dcache_nodeOut_a_bits_data = dcache_nodeOut_a_deq_bits_data ; 
    reg dcache_s1_valid ; 
    wire dcache_s1_valid_masked = dcache_s1_valid &~ dcache_io_cpu_s1_kill ; 
    wire dcache_s1_nack ; 
    wire dcache_s1_valid_not_nacked = dcache_s1_valid &~ dcache_s1_nack ; 
    wire dcache_s0_clk_en =(~ dcache_metaArb_grant_7 | dcache_io_cpu_req_valid )&~( dcache_metaArb_io_in_2_valid | dcache_metaArb_io_in_3_valid ); 
    wire[31:0] dcache_s0_tlb_req_vaddr = dcache_s0_req_addr ; 
    wire[4:0] dcache_s0_tlb_req_cmd = dcache_s0_req_cmd ; 
    wire[1:0] dcache_s0_tlb_req_size = dcache_s0_req_size ; 
    wire[1:0] dcache_s0_tlb_req_prv = dcache_s0_req_dprv ; 
    wire dcache_s0_tlb_req_v = dcache_s0_req_dv ; 
    wire dcache_s0_tlb_req_passthrough = dcache_s0_req_phys ; 
  assign  dcache_s0_req_addr ={ dcache_metaArb_io_in_2_valid | dcache_metaArb_io_in_3_valid  ? { dcache__metaArb_io_in_5_bits_addr_T , dcache_s2_vaddr [13:6]}: dcache_io_cpu_req_bits_addr [31:6], dcache_io_cpu_req_bits_addr [5:0]}; 
  assign  dcache_s0_req_phys =~ dcache_metaArb_grant_7 | dcache_io_cpu_req_bits_phys ; 
    wire[31:0] dcache_s1_vaddr = dcache_s1_req_addr ; reg[6:0] dcache_s1_req_tag ; 
    wire[1:0] dcache_s1_mask_xwr_size = dcache_s1_req_size ; 
    reg dcache_s1_req_signed ; 
    reg dcache_s1_req_dv ; 
    reg dcache_s1_req_phys ; 
    reg dcache_s1_req_no_xcpt ; 
    reg dcache_s1_tlb_req_passthrough ; 
    reg dcache_s1_tlb_req_v ; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_1 = dcache_s1_req_cmd ==5'h0; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_2 = dcache_s1_req_cmd ==5'h10; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_3 = dcache_s1_req_cmd ==5'h6; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_29 = dcache_s1_req_cmd ==5'h7; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_31 = dcache_s1_req_cmd ==5'h4; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_32 = dcache_s1_req_cmd ==5'h9; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_33 = dcache_s1_req_cmd ==5'hA; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_34 = dcache_s1_req_cmd ==5'hB; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_38 = dcache_s1_req_cmd ==5'h8; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_39 = dcache_s1_req_cmd ==5'hC; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_40 = dcache_s1_req_cmd ==5'hD; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_41 = dcache_s1_req_cmd ==5'hE; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_42 = dcache_s1_req_cmd ==5'hF; 
    wire dcache_s1_read = dcache__io_cpu_perf_canAcceptLoadThenLoad_T_1 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_2 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_3 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_29 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_31 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_32 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_33 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_34 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_38 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_39 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_40 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_41 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_42 ; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_26 = dcache_s1_req_cmd ==5'h1; 
    wire dcache__io_cpu_perf_canAcceptLoadThenLoad_T_51 = dcache_s1_req_cmd ==5'h11; 
    wire dcache_s1_write = dcache__io_cpu_perf_canAcceptLoadThenLoad_T_26 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_51 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_29 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_31 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_32 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_33 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_34 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_38 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_39 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_40 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_41 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_42 ; 
    wire dcache_s1_readwrite = dcache_s1_read | dcache_s1_write ; 
    wire dcache_s1_sfence = dcache_s1_req_cmd ==5'h14| dcache_s1_req_cmd ==5'h15| dcache_s1_req_cmd ==5'h16; 
    wire dcache_s1_flush_line = dcache_s1_req_cmd ==5'h5& dcache_s1_req_size [0]; 
    reg dcache_s1_flush_valid ; 
    reg dcache_cached_grant_wait ; reg[1:0] dcache_refill_way ; 
    wire dcache__io_cpu_req_ready_T_4 =~ dcache_cached_grant_wait &~ dcache_s1_nack ; 
    reg dcache_uncachedInFlight_0 ; reg[31:0] dcache_uncachedReqs_0_addr ; 
    wire[31:0] dcache_uncachedResp_addr = dcache_uncachedReqs_0_addr ; reg[6:0] dcache_uncachedReqs_0_tag ; 
    wire[6:0] dcache_uncachedResp_tag = dcache_uncachedReqs_0_tag ; reg[4:0] dcache_uncachedReqs_0_cmd ; 
    wire[4:0] dcache_uncachedResp_cmd = dcache_uncachedReqs_0_cmd ; reg[1:0] dcache_uncachedReqs_0_size ; 
    wire[1:0] dcache_uncachedResp_size = dcache_uncachedReqs_0_size ; 
    reg dcache_uncachedReqs_0_signed ; 
    wire dcache_uncachedResp_signed = dcache_uncachedReqs_0_signed ; reg[1:0] dcache_uncachedReqs_0_dprv ; 
    wire[1:0] dcache_uncachedResp_dprv = dcache_uncachedReqs_0_dprv ; 
    reg dcache_uncachedReqs_0_dv ; 
    wire dcache_uncachedResp_dv = dcache_uncachedReqs_0_dv ; 
    reg dcache_uncachedReqs_0_phys ; 
    wire dcache_uncachedResp_phys = dcache_uncachedReqs_0_phys ; 
    reg dcache_uncachedReqs_0_no_alloc ; 
    wire dcache_uncachedResp_no_alloc = dcache_uncachedReqs_0_no_alloc ; 
    reg dcache_uncachedReqs_0_no_xcpt ; 
    wire dcache_uncachedResp_no_xcpt = dcache_uncachedReqs_0_no_xcpt ; reg[31:0] dcache_uncachedReqs_0_data ; 
    wire[31:0] dcache_uncachedResp_data = dcache_uncachedReqs_0_data ; reg[3:0] dcache_uncachedReqs_0_mask ; 
    wire[3:0] dcache_uncachedResp_mask = dcache_uncachedReqs_0_mask ; 
    wire dcache__pstore_drain_opportunistic_T = dcache_io_cpu_req_bits_cmd ==5'h0; 
    wire dcache__pstore_drain_opportunistic_T_1 = dcache_io_cpu_req_bits_cmd ==5'h10; 
    wire dcache__pstore_drain_opportunistic_T_2 = dcache_io_cpu_req_bits_cmd ==5'h6; 
    wire dcache__pstore_drain_opportunistic_T_28 = dcache_io_cpu_req_bits_cmd ==5'h7; 
    wire dcache__pstore_drain_opportunistic_T_30 = dcache_io_cpu_req_bits_cmd ==5'h4; 
    wire dcache__pstore_drain_opportunistic_T_31 = dcache_io_cpu_req_bits_cmd ==5'h9; 
    wire dcache__pstore_drain_opportunistic_T_32 = dcache_io_cpu_req_bits_cmd ==5'hA; 
    wire dcache__pstore_drain_opportunistic_T_33 = dcache_io_cpu_req_bits_cmd ==5'hB; 
    wire dcache__pstore_drain_opportunistic_T_37 = dcache_io_cpu_req_bits_cmd ==5'h8; 
    wire dcache__pstore_drain_opportunistic_T_38 = dcache_io_cpu_req_bits_cmd ==5'hC; 
    wire dcache__pstore_drain_opportunistic_T_39 = dcache_io_cpu_req_bits_cmd ==5'hD; 
    wire dcache__pstore_drain_opportunistic_T_40 = dcache_io_cpu_req_bits_cmd ==5'hE; 
    wire dcache__pstore_drain_opportunistic_T_41 = dcache_io_cpu_req_bits_cmd ==5'hF; 
    wire dcache_s0_read = dcache__pstore_drain_opportunistic_T | dcache__pstore_drain_opportunistic_T_1 | dcache__pstore_drain_opportunistic_T_2 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 ; 
    wire dcache__pstore_drain_opportunistic_T_25 = dcache_io_cpu_req_bits_cmd ==5'h1; 
    wire dcache__pstore_drain_opportunistic_res_T_1 = dcache_io_cpu_req_bits_cmd ==5'h3; 
    wire dcache_dataArb_io_in_3_valid_res =~( dcache__pstore_drain_opportunistic_T_25 | dcache__pstore_drain_opportunistic_res_T_1 ); 
    wire dcache__pstore_drain_opportunistic_T_50 = dcache_io_cpu_req_bits_cmd ==5'h11; 
  assign  dcache_dataArb_io_in_3_valid = dcache_io_cpu_req_valid & dcache_dataArb_io_in_3_valid_res ; 
  assign  dcache__metaArb_io_in_5_bits_addr_T = dcache_io_cpu_req_bits_addr [31:14]; 
  assign  dcache_dataArb_io_in_3_bits_addr = dcache_io_cpu_req_bits_addr [13:0]; 
    reg dcache_s1_did_read ; 
    wire dcache_s2_data_word_en = dcache_s1_did_read ; 
    wire dcache__GEN_47 =~ dcache_metaArb_grant_7 |~ dcache_dataArb_grant_3 & dcache_s0_read ; 
    wire dcache_s1_cmd_uses_tlb = dcache_s1_readwrite | dcache_s1_flush_line | dcache_s1_req_cmd ==5'h17; 
    wire dcache_tlb_invalidate_refill = dcache_s1_valid &~ dcache_io_cpu_s1_kill & dcache_s1_sfence ; 
    wire[31:0] dcache_s1_paddr ={ dcache_tlb_ppn , dcache_s1_req_addr [11:0]}; 
    wire dcache_s1_hit_way = dcache_s1_paddr [31]& dcache_s1_paddr <32'h80004000; 
    wire[1:0] dcache_s1_hit_state_state ={2{ dcache_s1_hit_way }}; 
    wire[15:0] dcache_tl_d_data_encoded_lo = dcache_nodeOut_d_bits_data [15:0]; 
    wire[15:0] dcache_tl_d_data_encoded_lo_1 = dcache_nodeOut_d_bits_data [15:0]; 
    wire[15:0] dcache_tl_d_data_encoded_hi = dcache_nodeOut_d_bits_data [31:16]; 
    wire[15:0] dcache_tl_d_data_encoded_hi_1 = dcache_nodeOut_d_bits_data [31:16]; 
    wire[31:0] dcache_s1_all_data_ways_1 = dcache_tl_d_data_encoded ; 
    wire[31:0] dcache_s2_data_s1_way_words_0_0 = dcache_s1_all_data_ways_0 ; 
    wire[31:0] dcache_s2_data_s1_way_words_1_0 = dcache_s1_all_data_ways_1 ; 
    wire dcache_s1_mask_xwr_upper = dcache_s1_req_addr [0]|(| dcache_s1_mask_xwr_size ); 
    wire dcache_s1_mask_xwr_lower =~( dcache_s1_req_addr [0]); 
    wire[1:0] dcache__s1_mask_xwr_T ={ dcache_s1_mask_xwr_upper , dcache_s1_mask_xwr_lower }; 
    wire[1:0] dcache_s1_mask_xwr_upper_1 =( dcache_s1_req_addr [1] ?  dcache__s1_mask_xwr_T :2'h0)|{2{ dcache_s1_mask_xwr_size [1]}}; 
    wire[1:0] dcache_s1_mask_xwr_lower_1 = dcache_s1_req_addr [1] ? 2'h0: dcache__s1_mask_xwr_T ; 
    wire[3:0] dcache_s1_mask_xwr ={ dcache_s1_mask_xwr_upper_1 , dcache_s1_mask_xwr_lower_1 }; 
    wire[3:0] dcache_s1_mask = dcache__io_cpu_perf_canAcceptLoadThenLoad_T_51  ?  dcache_io_cpu_s1_data_mask : dcache_s1_mask_xwr ; 
    reg dcache_s2_valid ; 
    wire[1:0] dcache_s2_valid_no_xcpt_lo_lo ={ dcache__io_cpu_s2_xcpt_ae_ld_output , dcache__io_cpu_s2_xcpt_ae_st_output }; 
    wire[3:0] dcache_s2_valid_no_xcpt_lo ={2'h0, dcache_s2_valid_no_xcpt_lo_lo }; 
    wire[1:0] dcache_s2_valid_no_xcpt_hi_lo ={ dcache__io_cpu_s2_xcpt_pf_ld_output , dcache__io_cpu_s2_xcpt_pf_st_output }; 
    wire[1:0] dcache_s2_valid_no_xcpt_hi_hi ={ dcache__io_cpu_s2_xcpt_ma_ld_output , dcache__io_cpu_s2_xcpt_ma_st_output }; 
    wire[3:0] dcache_s2_valid_no_xcpt_hi ={ dcache_s2_valid_no_xcpt_hi_hi , dcache_s2_valid_no_xcpt_hi_lo }; 
    wire dcache_s2_valid_no_xcpt = dcache_s2_valid &{ dcache_s2_valid_no_xcpt_hi , dcache_s2_valid_no_xcpt_lo }==8'h0; 
    reg dcache_s2_not_nacked_in_s1 ; 
    wire dcache_s2_valid_not_nacked_in_s1 = dcache_s2_valid & dcache_s2_not_nacked_in_s1 ; 
    wire dcache_s2_valid_masked = dcache_s2_valid_no_xcpt & dcache_s2_not_nacked_in_s1 ; 
    wire dcache_s2_valid_not_killed = dcache_s2_valid_masked ; reg[31:0] dcache_s2_req_addr ; 
    wire[31:0] dcache_get_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_put_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_putpartial_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_1_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_2_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_3_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_4_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_5_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_6_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_7_address = dcache_s2_req_addr ; 
    wire[31:0] dcache_atomics_a_8_address = dcache_s2_req_addr ; reg[6:0] dcache_s2_req_tag ; reg[4:0] dcache_s2_req_cmd ; reg[1:0] dcache_s2_req_size ; 
    wire[1:0] dcache_size = dcache_s2_req_size ; 
    reg dcache_s2_req_signed ; reg[1:0] dcache_s2_req_dprv ; 
    reg dcache_s2_req_dv ; 
    reg dcache_s2_req_phys ; 
    reg dcache_s2_req_no_alloc ; 
    reg dcache_s2_req_no_xcpt ; reg[31:0] dcache_s2_req_data ; reg[3:0] dcache_s2_req_mask ; 
    wire dcache__s2_cmd_flush_line_T = dcache_s2_req_cmd ==5'h5; 
    wire dcache_s2_cmd_flush_all = dcache__s2_cmd_flush_line_T &~( dcache_s2_req_size [0]); 
    wire dcache_s2_cmd_flush_line = dcache__s2_cmd_flush_line_T & dcache_s2_req_size [0]; reg[31:0] dcache_s2_tlb_xcpt_paddr ; reg[31:0] dcache_s2_tlb_xcpt_gpa ; 
    reg dcache_s2_tlb_xcpt_pf_ld ; 
    reg dcache_s2_tlb_xcpt_pf_st ; 
    reg dcache_s2_tlb_xcpt_pf_inst ; 
    reg dcache_s2_tlb_xcpt_ae_ld ; 
    reg dcache_s2_tlb_xcpt_ae_st ; 
    reg dcache_s2_tlb_xcpt_ae_inst ; 
    reg dcache_s2_tlb_xcpt_ma_ld ; 
    reg dcache_s2_tlb_xcpt_ma_st ; 
    reg dcache_s2_tlb_xcpt_cacheable ; 
    reg dcache_s2_tlb_xcpt_must_alloc ; 
    reg dcache_s2_tlb_xcpt_prefetchable ; reg[31:0] dcache_s2_pma_paddr ; reg[31:0] dcache_s2_pma_gpa ; 
    reg dcache_s2_pma_pf_ld ; 
    reg dcache_s2_pma_pf_st ; 
    reg dcache_s2_pma_pf_inst ; 
    reg dcache_s2_pma_ae_ld ; 
    reg dcache_s2_pma_ae_st ; 
    reg dcache_s2_pma_ae_inst ; 
    reg dcache_s2_pma_ma_ld ; 
    reg dcache_s2_pma_ma_st ; 
    reg dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_bufferable = dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_modifiable = dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_readalloc = dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_writealloc = dcache_s2_pma_cacheable ; 
    reg dcache_s2_pma_must_alloc ; 
    reg dcache_s2_pma_prefetchable ; reg[31:0] dcache_s2_uncached_resp_addr ; 
    wire dcache_s1_meta_clk_en = dcache_s1_valid_not_nacked | dcache_s1_flush_valid ; reg[31:0] dcache_s2_vaddr_r ; 
  assign  dcache_s2_vaddr ={ dcache_s2_vaddr_r [31:14], dcache_s2_req_addr [13:0]}; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_48 = dcache_s2_req_cmd ==5'h6; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_26 = dcache_s2_req_cmd ==5'h7; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_28 = dcache_s2_req_cmd ==5'h4; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_29 = dcache_s2_req_cmd ==5'h9; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_30 = dcache_s2_req_cmd ==5'hA; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_31 = dcache_s2_req_cmd ==5'hB; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_35 = dcache_s2_req_cmd ==5'h8; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_36 = dcache_s2_req_cmd ==5'hC; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_37 = dcache_s2_req_cmd ==5'hD; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_38 = dcache_s2_req_cmd ==5'hE; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_39 = dcache_s2_req_cmd ==5'hF; 
    wire dcache_s2_read = dcache_s2_req_cmd ==5'h0| dcache_s2_req_cmd ==5'h10| dcache__metaArb_io_in_3_bits_data_c_cat_T_48 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 | dcache__metaArb_io_in_3_bits_data_c_cat_T_28 | dcache__metaArb_io_in_3_bits_data_c_cat_T_29 | dcache__metaArb_io_in_3_bits_data_c_cat_T_30 | dcache__metaArb_io_in_3_bits_data_c_cat_T_31 | dcache__metaArb_io_in_3_bits_data_c_cat_T_35 | dcache__metaArb_io_in_3_bits_data_c_cat_T_36 | dcache__metaArb_io_in_3_bits_data_c_cat_T_37 | dcache__metaArb_io_in_3_bits_data_c_cat_T_38 | dcache__metaArb_io_in_3_bits_data_c_cat_T_39 ; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_23 = dcache_s2_req_cmd ==5'h1; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_24 = dcache_s2_req_cmd ==5'h11; 
    wire dcache_s2_write = dcache__metaArb_io_in_3_bits_data_c_cat_T_23 | dcache__metaArb_io_in_3_bits_data_c_cat_T_24 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 | dcache__metaArb_io_in_3_bits_data_c_cat_T_28 | dcache__metaArb_io_in_3_bits_data_c_cat_T_29 | dcache__metaArb_io_in_3_bits_data_c_cat_T_30 | dcache__metaArb_io_in_3_bits_data_c_cat_T_31 | dcache__metaArb_io_in_3_bits_data_c_cat_T_35 | dcache__metaArb_io_in_3_bits_data_c_cat_T_36 | dcache__metaArb_io_in_3_bits_data_c_cat_T_37 | dcache__metaArb_io_in_3_bits_data_c_cat_T_38 | dcache__metaArb_io_in_3_bits_data_c_cat_T_39 ; 
    wire dcache_s2_readwrite = dcache_s2_read | dcache_s2_write ; 
    reg dcache_s2_flush_valid_pre_tag_ecc ; 
    wire dcache_s2_flush_valid = dcache_s2_flush_valid_pre_tag_ecc ; 
    wire dcache_s2_data_en = dcache_s1_valid | dcache__io_cpu_replay_next_output ; 
    wire dcache_s2_data_s1_word_en = dcache__io_cpu_replay_next_output | dcache_s2_data_word_en ; reg[31:0] dcache_s2_data ; 
    reg dcache_s2_probe_way ; 
    wire dcache_releaseWay = dcache_s2_probe_way ; reg[1:0] dcache_s2_probe_state_state ; 
    reg dcache_s2_hit_way ; reg[1:0] dcache_s2_hit_state_state ; 
    wire dcache_s2_hit_valid =| dcache_s2_hit_state_state ; 
    wire dcache__metaArb_io_in_3_bits_data_c_cat_T_46 = dcache_s2_req_cmd ==5'h3; 
    wire[1:0] dcache_c ={ dcache__metaArb_io_in_3_bits_data_c_cat_T_23 | dcache__metaArb_io_in_3_bits_data_c_cat_T_24 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 | dcache__metaArb_io_in_3_bits_data_c_cat_T_28 | dcache__metaArb_io_in_3_bits_data_c_cat_T_29 | dcache__metaArb_io_in_3_bits_data_c_cat_T_30 | dcache__metaArb_io_in_3_bits_data_c_cat_T_31 | dcache__metaArb_io_in_3_bits_data_c_cat_T_35 | dcache__metaArb_io_in_3_bits_data_c_cat_T_36 | dcache__metaArb_io_in_3_bits_data_c_cat_T_37 | dcache__metaArb_io_in_3_bits_data_c_cat_T_38 | dcache__metaArb_io_in_3_bits_data_c_cat_T_39 , dcache__metaArb_io_in_3_bits_data_c_cat_T_23 | dcache__metaArb_io_in_3_bits_data_c_cat_T_24 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 | dcache__metaArb_io_in_3_bits_data_c_cat_T_28 | dcache__metaArb_io_in_3_bits_data_c_cat_T_29 | dcache__metaArb_io_in_3_bits_data_c_cat_T_30 | dcache__metaArb_io_in_3_bits_data_c_cat_T_31 | dcache__metaArb_io_in_3_bits_data_c_cat_T_35 | dcache__metaArb_io_in_3_bits_data_c_cat_T_36 | dcache__metaArb_io_in_3_bits_data_c_cat_T_37 | dcache__metaArb_io_in_3_bits_data_c_cat_T_38 | dcache__metaArb_io_in_3_bits_data_c_cat_T_39 | dcache__metaArb_io_in_3_bits_data_c_cat_T_46 | dcache__metaArb_io_in_3_bits_data_c_cat_T_48 }; 
    wire[3:0] dcache__GEN_48 ={ dcache_c , dcache_s2_hit_state_state }; 
    wire dcache_s2_hit = dcache__GEN_48 ==4'h3| dcache__GEN_48 ==4'h2| dcache__GEN_48 ==4'h1| dcache__GEN_48 ==4'h7| dcache__GEN_48 ==4'h6|(& dcache__GEN_48 )| dcache__GEN_48 ==4'hE; reg[1:0] dcache_casez_tmp ; 
    wire[1:0] dcache__GEN_49 ={1'h0, dcache__GEN_48 ==4'hC}; 
  always @(*)
         begin 
             casez ( dcache__GEN_48 )
              4 'b0000: 
                  dcache_casez_tmp  =2'h0;
              4 'b0001: 
                  dcache_casez_tmp  =2'h1;
              4 'b0010: 
                  dcache_casez_tmp  =2'h2;
              4 'b0011: 
                  dcache_casez_tmp  =2'h3;
              4 'b0100: 
                  dcache_casez_tmp  =2'h1;
              4 'b0101: 
                  dcache_casez_tmp  =2'h2;
              4 'b0110: 
                  dcache_casez_tmp  =2'h2;
              4 'b0111: 
                  dcache_casez_tmp  =2'h3;
              4 'b1000: 
                  dcache_casez_tmp  = dcache__GEN_49 ;
              4 'b1001: 
                  dcache_casez_tmp  = dcache__GEN_49 ;
              4 'b1010: 
                  dcache_casez_tmp  = dcache__GEN_49 ;
              4 'b1011: 
                  dcache_casez_tmp  = dcache__GEN_49 ;
              4 'b1100: 
                  dcache_casez_tmp  = dcache__GEN_49 ;
              4 'b1101: 
                  dcache_casez_tmp  =2'h2;
              4 'b1110: 
                  dcache_casez_tmp  =2'h3;
              default : 
                  dcache_casez_tmp  =2'h3;endcase
         end
    wire[1:0] dcache_s2_grow_param = dcache_casez_tmp ; 
    wire[1:0] dcache_s2_new_hit_state_state = dcache_s2_grow_param ; 
    wire[1:0] dcache_metaArb_io_in_2_bits_data_meta_coh_state = dcache_s2_new_hit_state_state ; 
    wire[15:0] dcache_s2_data_corrected_lo = dcache_s2_data [15:0]; 
    wire[15:0] dcache_s2_data_uncorrected_lo = dcache_s2_data [15:0]; 
    wire[15:0] dcache_s2_data_corrected_hi = dcache_s2_data [31:16]; 
    wire[15:0] dcache_s2_data_uncorrected_hi = dcache_s2_data [31:16]; 
    wire[31:0] dcache_s2_data_corrected ={ dcache_s2_data_corrected_hi , dcache_s2_data_corrected_lo }; 
    wire[31:0] dcache_s2_data_word_corrected = dcache_s2_data_corrected ; 
    wire[31:0] dcache_s2_data_uncorrected ={ dcache_s2_data_uncorrected_hi , dcache_s2_data_uncorrected_lo }; 
    wire[31:0] dcache_s2_data_word = dcache_s2_data_uncorrected ; 
    wire dcache_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = dcache_s2_valid_masked & dcache_s2_hit ; 
    wire dcache_s2_valid_hit_pre_data_ecc_and_waw = dcache_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & dcache_s2_readwrite ; 
    wire dcache_s2_valid_hit_pre_data_ecc = dcache_s2_valid_hit_pre_data_ecc_and_waw ; 
    wire dcache_s2_valid_flush_line = dcache_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & dcache_s2_cmd_flush_line ; 
    wire dcache_s2_valid_hit = dcache_s2_valid_hit_pre_data_ecc ; 
    wire dcache_s2_valid_miss = dcache_s2_valid_masked & dcache_s2_readwrite &~ dcache_s2_hit ; 
    wire dcache_s2_uncached =~ dcache_s2_pma_cacheable | dcache_s2_req_no_alloc &~ dcache_s2_pma_must_alloc &~ dcache_s2_hit_valid ; 
    wire dcache_s2_valid_cached_miss = dcache_s2_valid_miss &~ dcache_s2_uncached &~ dcache_uncachedInFlight_0 ; 
    wire dcache_s2_valid_uncached_pending = dcache_s2_valid_miss & dcache_s2_uncached &~ dcache_uncachedInFlight_0 ; 
    wire[1:0] dcache_s2_victim_or_hit_way = dcache_s2_hit_valid  ? {1'h0, dcache_s2_hit_way }:2'h1; 
    wire[17:0] dcache_s2_victim_tag = dcache_s2_valid_flush_line  ?  dcache_s2_req_addr [31:14]:18'h0; 
    wire[1:0] dcache_s2_victim_state_state = dcache_s2_hit_valid  ?  dcache_s2_hit_state_state :2'h0; 
    wire dcache__GEN_50 = dcache_s2_probe_state_state ==2'h1; 
    wire dcache_s2_prb_ack_data =& dcache_s2_probe_state_state ; 
    wire dcache__GEN_51 =(& dcache_s2_probe_state_state )| dcache_s2_probe_state_state ==2'h2; 
    wire[2:0] dcache_s2_report_param = dcache__GEN_51  ? 3'h3: dcache__GEN_50  ? 3'h4: dcache_s2_probe_state_state ==2'h0 ? 3'h5:3'h0; 
    wire[2:0] dcache_cleanReleaseMessage_param = dcache_s2_report_param ; 
    wire[2:0] dcache_dirtyReleaseMessage_param = dcache_s2_report_param ; 
    wire[1:0] dcache_probeNewCoh_state = dcache__GEN_51  ? 2'h2:{1'h0, dcache__GEN_50 }; 
    wire[1:0] dcache_newCoh_state = dcache_probeNewCoh_state ; 
    wire[2:0] dcache_s2_shrink_param =(& dcache_s2_victim_state_state )| dcache_s2_victim_state_state ==2'h2 ? 3'h1: dcache_s2_victim_state_state ==2'h1 ? 3'h2: dcache_s2_victim_state_state ==2'h0 ? 3'h5:3'h0; 
    wire dcache_s2_victim_dirty =& dcache_s2_victim_state_state ; 
    wire dcache_s2_update_meta = dcache_s2_hit_state_state != dcache_s2_new_hit_state_state ; 
    wire dcache_s2_dont_nack_uncached = dcache_s2_valid_uncached_pending & dcache_tl_out_a_ready ; 
    wire dcache_s2_dont_nack_misc = dcache_s2_valid_masked & dcache_s2_req_cmd ==5'h17; 
    wire dcache__io_cpu_s2_nack_output = dcache_s2_valid_no_xcpt &~ dcache_s2_dont_nack_uncached &~ dcache_s2_dont_nack_misc &~ dcache_s2_valid_hit ; 
  assign  dcache_metaArb_io_in_2_valid = dcache_s2_valid_hit_pre_data_ecc_and_waw & dcache_s2_update_meta ; 
    wire[17:0] dcache_metaArb_io_in_2_bits_data_meta_tag = dcache_s2_req_addr [31:14]; 
    wire[17:0] dcache_metaArb_io_in_3_bits_data_meta_1_tag = dcache_s2_req_addr [31:14]; reg[6:0] dcache_lrscCount ; 
    wire dcache_lrscValid =|( dcache_lrscCount [6:2]); 
    wire dcache_lrscBackingOff =(| dcache_lrscCount )&~ dcache_lrscValid ; reg[25:0] dcache_lrscAddr ; 
    wire dcache_lrscAddrMatch = dcache_lrscAddr == dcache_s2_req_addr [31:6]; 
    reg dcache_s2_correct_REG ; reg[4:0] dcache_pstore1_cmd ; reg[31:0] dcache_pstore1_addr ; reg[31:0] dcache_pstore1_data ; 
    wire[31:0] dcache_put_data = dcache_pstore1_data ; 
    wire[31:0] dcache_putpartial_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_1_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_2_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_3_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_4_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_5_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_6_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_7_data = dcache_pstore1_data ; 
    wire[31:0] dcache_atomics_a_8_data = dcache_pstore1_data ; 
    reg dcache_pstore1_way ; reg[3:0] dcache_pstore1_mask ; 
    wire[3:0] dcache_pstore2_storegen_mask_mergedMask = dcache_pstore1_mask ; 
    reg dcache_pstore1_rmw_r ; 
    wire dcache_pstore1_rmw = dcache_pstore1_rmw_r ; 
    wire dcache__pstore1_held_T = dcache_s2_valid_hit & dcache_s2_write ; 
    reg dcache_pstore2_valid ; 
    wire dcache_pstore_drain_opportunistic_res =~( dcache__pstore_drain_opportunistic_T_25 | dcache__pstore_drain_opportunistic_res_T_1 ); 
    wire dcache_pstore_drain_opportunistic =~( dcache_io_cpu_req_valid & dcache_pstore_drain_opportunistic_res ); 
    reg dcache_pstore_drain_on_miss_REG ; 
    wire dcache_pstore_drain_on_miss = dcache_pstore_drain_on_miss_REG ; 
    reg dcache_pstore1_held ; 
    wire dcache_pstore1_valid_likely = dcache_s2_valid & dcache_s2_write | dcache_pstore1_held ; 
    wire dcache_pstore1_valid = dcache__pstore1_held_T | dcache_pstore1_held ; 
    wire dcache_any_pstore_valid = dcache_pstore1_held | dcache_pstore2_valid ; 
    wire dcache_pstore_drain_structural = dcache_pstore1_valid_likely & dcache_pstore2_valid &( dcache_s1_valid & dcache_s1_write | dcache_pstore1_rmw ); 
    wire dcache__dataArb_io_in_0_valid_T_2 = dcache_s2_valid_hit_pre_data_ecc & dcache_s2_write ; 
    wire dcache__dataArb_io_in_0_valid_T_9 = dcache_pstore_drain_opportunistic | dcache_pstore_drain_on_miss ; 
  assign  dcache_pstore_drain = dcache_pstore_drain_structural |(( dcache__dataArb_io_in_0_valid_T_2 | dcache_pstore1_held )&~ dcache_pstore1_rmw | dcache_pstore2_valid )& dcache__dataArb_io_in_0_valid_T_9 ; 
    wire dcache_advance_pstore1 = dcache_pstore1_valid & dcache_pstore2_valid == dcache_pstore_drain ; reg[31:0] dcache_pstore2_addr ; 
    reg dcache_pstore2_way ; reg[7:0] dcache_pstore2_storegen_data_r ; reg[7:0] dcache_pstore2_storegen_data_r_1 ; reg[7:0] dcache_pstore2_storegen_data_r_2 ; reg[7:0] dcache_pstore2_storegen_data_r_3 ; 
    wire[15:0] dcache_pstore2_storegen_data_lo ={ dcache_pstore2_storegen_data_r_1 , dcache_pstore2_storegen_data_r }; 
    wire[15:0] dcache_pstore2_storegen_data_hi ={ dcache_pstore2_storegen_data_r_3 , dcache_pstore2_storegen_data_r_2 }; 
    wire[31:0] dcache_pstore2_storegen_data ={ dcache_pstore2_storegen_data_hi , dcache_pstore2_storegen_data_lo }; reg[3:0] dcache_pstore2_storegen_mask ; 
  assign  dcache_dataArb_io_in_0_valid = dcache_pstore_drain_structural |(( dcache__dataArb_io_in_0_valid_T_2 | dcache_pstore1_held )&~ dcache_pstore1_rmw | dcache_pstore2_valid )& dcache__dataArb_io_in_0_valid_T_9 ; 
  assign  dcache__dataArb_io_in_0_bits_wordMask_wordMask_T = dcache_pstore2_valid  ?  dcache_pstore2_addr [13:0]: dcache_pstore1_addr [13:0]; 
    wire[31:0] dcache__dataArb_io_in_0_bits_wdata_T = dcache_pstore2_valid  ?  dcache_pstore2_storegen_data : dcache_pstore1_data ; 
    wire[15:0] dcache_dataArb_io_in_0_bits_wdata_lo = dcache__dataArb_io_in_0_bits_wdata_T [15:0]; 
    wire[15:0] dcache_dataArb_io_in_0_bits_wdata_hi = dcache__dataArb_io_in_0_bits_wdata_T [31:16]; 
    wire[1:0] dcache_dataArb_io_in_0_bits_eccMask_hi ; 
    wire[1:0] dcache_dataArb_io_in_0_bits_eccMask_lo ; 
    wire dcache_dataArb_io_in_0_bits_wordMask_eccMask =(| dcache_dataArb_io_in_0_bits_eccMask_lo )| dcache_dataArb_io_in_0_bits_eccMask_hi [0]| dcache_dataArb_io_in_0_bits_eccMask_hi [1]; 
    wire[3:0] dcache__dataArb_io_in_0_bits_eccMask_T = dcache_pstore2_valid  ?  dcache_pstore2_storegen_mask : dcache_pstore1_mask ; 
  assign  dcache_dataArb_io_in_0_bits_eccMask_lo = dcache__dataArb_io_in_0_bits_eccMask_T [1:0]; 
  assign  dcache_dataArb_io_in_0_bits_eccMask_hi = dcache__dataArb_io_in_0_bits_eccMask_T [3:2]; 
  assign  dcache_dataArb_io_in_1_bits_eccMask ={ dcache_dataArb_io_in_0_bits_eccMask_hi , dcache_dataArb_io_in_0_bits_eccMask_lo }; 
    wire[1:0] dcache_s1_hazard_lo = dcache_pstore1_mask [1:0]; 
    wire[1:0] dcache_s1_hazard_lo_1 = dcache_s1_hazard_lo ; 
    wire[1:0] dcache_s1_hazard_hi = dcache_pstore1_mask [3:2]; 
    wire[1:0] dcache_s1_hazard_hi_1 = dcache_s1_hazard_hi ; 
    wire[1:0] dcache_s1_hazard_lo_2 = dcache_s1_mask_xwr [1:0]; 
    wire[1:0] dcache_s1_hazard_lo_6 = dcache_s1_mask_xwr [1:0]; 
    wire[1:0] dcache_s1_hazard_lo_3 = dcache_s1_hazard_lo_2 ; 
    wire[1:0] dcache_s1_hazard_hi_2 = dcache_s1_mask_xwr [3:2]; 
    wire[1:0] dcache_s1_hazard_hi_6 = dcache_s1_mask_xwr [3:2]; 
    wire[1:0] dcache_s1_hazard_hi_3 = dcache_s1_hazard_hi_2 ; 
    wire[1:0] dcache_s1_hazard_lo_4 = dcache_pstore2_storegen_mask [1:0]; 
    wire[1:0] dcache_s1_hazard_lo_5 = dcache_s1_hazard_lo_4 ; 
    wire[1:0] dcache_s1_hazard_hi_4 = dcache_pstore2_storegen_mask [3:2]; 
    wire[1:0] dcache_s1_hazard_hi_5 = dcache_s1_hazard_hi_4 ; 
    wire[1:0] dcache_s1_hazard_lo_7 = dcache_s1_hazard_lo_6 ; 
    wire[1:0] dcache_s1_hazard_hi_7 = dcache_s1_hazard_hi_6 ; 
    wire dcache_s1_hazard = dcache_pstore1_valid_likely & dcache_pstore1_addr [13:2]== dcache_s1_vaddr [13:2]&( dcache_s1_write  ? (|({ dcache_s1_hazard_hi_1 , dcache_s1_hazard_lo_1 }&{ dcache_s1_hazard_hi_3 , dcache_s1_hazard_lo_3 })):(|( dcache_pstore1_mask & dcache_s1_mask_xwr )))| dcache_pstore2_valid & dcache_pstore2_addr [13:2]== dcache_s1_vaddr [13:2]&( dcache_s1_write  ? (|({ dcache_s1_hazard_hi_5 , dcache_s1_hazard_lo_5 }&{ dcache_s1_hazard_hi_7 , dcache_s1_hazard_lo_7 })):(|( dcache_pstore2_storegen_mask & dcache_s1_mask_xwr ))); 
    wire dcache_s1_raw_hazard = dcache_s1_read & dcache_s1_hazard ; 
  assign  dcache_s1_nack = dcache_s1_valid & dcache_s1_raw_hazard | dcache__io_cpu_s2_nack_output | dcache_metaArb_io_in_2_valid ; 
    reg dcache_io_cpu_s2_nack_cause_raw_REG ; 
    wire[31:0] dcache__GEN_52 ={ dcache_s2_req_addr [31:6],6'h0}; 
    wire[31:0] dcache_acquire_address ; 
  assign  dcache_acquire_address = dcache__GEN_52 ; 
    wire[31:0] dcache_error_addr ; 
  assign  dcache_error_addr = dcache__GEN_52 ; 
    wire[18:0] dcache_a_mask ={15'h0, dcache_pstore1_mask }; 
    wire[5:0] dcache__GEN_53 ={ dcache_s2_req_addr [31:30], dcache_s2_req_addr [27], dcache_s2_req_addr [25], dcache_s2_req_addr [16],~( dcache_s2_req_addr [13])}; 
    wire[5:0] dcache__GEN_54 ={ dcache_s2_req_addr [31:30], dcache_s2_req_addr [27], dcache_s2_req_addr [25], dcache_s2_req_addr [16], dcache_s2_req_addr [13]}; 
    wire[4:0] dcache__GEN_55 ={ dcache_s2_req_addr [31:30], dcache_s2_req_addr [27],~( dcache_s2_req_addr [25]), dcache_s2_req_addr [16]}; 
    wire[2:0] dcache__GEN_56 ={ dcache_s2_req_addr [31:30],~( dcache_s2_req_addr [27])}; 
    wire[1:0] dcache__GEN_57 ={ dcache_s2_req_addr [31],~( dcache_s2_req_addr [30])}; 
    wire[4:0] dcache__GEN_58 ={ dcache_s2_req_addr [31:30]^2'h2, dcache_s2_req_addr [27], dcache_s2_req_addr [25], dcache_s2_req_addr [16]}; 
    wire dcache_get_legal =~(| dcache__GEN_53 )|~(| dcache__GEN_54 )|{ dcache_s2_req_addr [31:30], dcache_s2_req_addr [27], dcache_s2_req_addr [25],~( dcache_s2_req_addr [16])}==5'h0|~(| dcache__GEN_55 )|~(| dcache__GEN_56 )|~(| dcache__GEN_57 )|~(| dcache__GEN_58 ); 
    wire[3:0] dcache__GEN_59 ={2'h0, dcache_s2_req_size }; 
    wire[3:0] dcache_get_size ; 
  assign  dcache_get_size = dcache__GEN_59 ; 
    wire[3:0] dcache_put_size ; 
  assign  dcache_put_size = dcache__GEN_59 ; 
    wire[3:0] dcache_putpartial_size ; 
  assign  dcache_putpartial_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_size ; 
  assign  dcache_atomics_a_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_1_size ; 
  assign  dcache_atomics_a_1_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_2_size ; 
  assign  dcache_atomics_a_2_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_3_size ; 
  assign  dcache_atomics_a_3_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_4_size ; 
  assign  dcache_atomics_a_4_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_5_size ; 
  assign  dcache_atomics_a_5_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_6_size ; 
  assign  dcache_atomics_a_6_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_7_size ; 
  assign  dcache_atomics_a_7_size = dcache__GEN_59 ; 
    wire[3:0] dcache_atomics_a_8_size ; 
  assign  dcache_atomics_a_8_size = dcache__GEN_59 ; 
    wire dcache_get_a_mask_sizeOH_shiftAmount = dcache_s2_req_size [0]; 
    wire dcache_put_a_mask_sizeOH_shiftAmount = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_1 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_2 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_3 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_4 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_5 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_6 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_7 = dcache_s2_req_size [0]; 
    wire dcache_atomics_a_mask_sizeOH_shiftAmount_8 = dcache_s2_req_size [0]; 
    wire[1:0] dcache_get_a_mask_sizeOH ={ dcache_get_a_mask_sizeOH_shiftAmount ,1'h1}; 
    wire dcache_get_a_mask_size = dcache_get_a_mask_sizeOH [1]; 
    wire dcache_get_a_mask_bit = dcache_s2_req_addr [1]; 
    wire dcache_put_a_mask_bit = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_2 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_4 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_6 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_8 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_10 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_12 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_14 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_bit_16 = dcache_s2_req_addr [1]; 
    wire dcache_get_a_mask_eq_1 = dcache_get_a_mask_bit ; 
    wire dcache_get_a_mask_nbit =~ dcache_get_a_mask_bit ; 
    wire dcache_get_a_mask_eq = dcache_get_a_mask_nbit ; 
    wire dcache_get_a_mask_acc = dcache_s2_req_size [1]| dcache_get_a_mask_size & dcache_get_a_mask_eq ; 
    wire dcache_get_a_mask_acc_1 = dcache_s2_req_size [1]| dcache_get_a_mask_size & dcache_get_a_mask_eq_1 ; 
    wire dcache_get_a_mask_size_1 = dcache_get_a_mask_sizeOH [0]; 
    wire dcache_get_a_mask_bit_1 = dcache_s2_req_addr [0]; 
    wire dcache_put_a_mask_bit_1 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_1 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_3 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_5 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_7 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_9 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_11 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_13 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_15 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_bit_17 = dcache_s2_req_addr [0]; 
    wire dcache_get_a_mask_nbit_1 =~ dcache_get_a_mask_bit_1 ; 
    wire dcache_get_a_mask_eq_2 = dcache_get_a_mask_eq & dcache_get_a_mask_nbit_1 ; 
    wire dcache_get_a_mask_acc_2 = dcache_get_a_mask_acc | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_2 ; 
    wire dcache_get_a_mask_eq_3 = dcache_get_a_mask_eq & dcache_get_a_mask_bit_1 ; 
    wire dcache_get_a_mask_acc_3 = dcache_get_a_mask_acc | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_3 ; 
    wire dcache_get_a_mask_eq_4 = dcache_get_a_mask_eq_1 & dcache_get_a_mask_nbit_1 ; 
    wire dcache_get_a_mask_acc_4 = dcache_get_a_mask_acc_1 | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_4 ; 
    wire dcache_get_a_mask_eq_5 = dcache_get_a_mask_eq_1 & dcache_get_a_mask_bit_1 ; 
    wire dcache_get_a_mask_acc_5 = dcache_get_a_mask_acc_1 | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_5 ; 
    wire[1:0] dcache_get_a_mask_lo ={ dcache_get_a_mask_acc_3 , dcache_get_a_mask_acc_2 }; 
    wire[1:0] dcache_get_a_mask_hi ={ dcache_get_a_mask_acc_5 , dcache_get_a_mask_acc_4 }; 
    wire[3:0] dcache_get_mask ={ dcache_get_a_mask_hi , dcache_get_a_mask_lo }; 
    wire dcache_put_legal =~(| dcache__GEN_53 )|~(| dcache__GEN_54 )|~(| dcache__GEN_55 )|~(| dcache__GEN_56 )|~(| dcache__GEN_58 )|~(| dcache__GEN_57 ); 
    wire[1:0] dcache_put_a_mask_sizeOH ={ dcache_put_a_mask_sizeOH_shiftAmount ,1'h1}; 
    wire dcache_put_a_mask_size = dcache_put_a_mask_sizeOH [1]; 
    wire dcache_put_a_mask_eq_1 = dcache_put_a_mask_bit ; 
    wire dcache_put_a_mask_nbit =~ dcache_put_a_mask_bit ; 
    wire dcache_put_a_mask_eq = dcache_put_a_mask_nbit ; 
    wire dcache_put_a_mask_acc = dcache_s2_req_size [1]| dcache_put_a_mask_size & dcache_put_a_mask_eq ; 
    wire dcache_put_a_mask_acc_1 = dcache_s2_req_size [1]| dcache_put_a_mask_size & dcache_put_a_mask_eq_1 ; 
    wire dcache_put_a_mask_size_1 = dcache_put_a_mask_sizeOH [0]; 
    wire dcache_put_a_mask_nbit_1 =~ dcache_put_a_mask_bit_1 ; 
    wire dcache_put_a_mask_eq_2 = dcache_put_a_mask_eq & dcache_put_a_mask_nbit_1 ; 
    wire dcache_put_a_mask_acc_2 = dcache_put_a_mask_acc | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_2 ; 
    wire dcache_put_a_mask_eq_3 = dcache_put_a_mask_eq & dcache_put_a_mask_bit_1 ; 
    wire dcache_put_a_mask_acc_3 = dcache_put_a_mask_acc | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_3 ; 
    wire dcache_put_a_mask_eq_4 = dcache_put_a_mask_eq_1 & dcache_put_a_mask_nbit_1 ; 
    wire dcache_put_a_mask_acc_4 = dcache_put_a_mask_acc_1 | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_4 ; 
    wire dcache_put_a_mask_eq_5 = dcache_put_a_mask_eq_1 & dcache_put_a_mask_bit_1 ; 
    wire dcache_put_a_mask_acc_5 = dcache_put_a_mask_acc_1 | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_5 ; 
    wire[1:0] dcache_put_a_mask_lo ={ dcache_put_a_mask_acc_3 , dcache_put_a_mask_acc_2 }; 
    wire[1:0] dcache_put_a_mask_hi ={ dcache_put_a_mask_acc_5 , dcache_put_a_mask_acc_4 }; 
    wire[3:0] dcache_put_mask ={ dcache_put_a_mask_hi , dcache_put_a_mask_lo }; 
    wire dcache_putpartial_legal =~(| dcache__GEN_53 )|~(| dcache__GEN_54 )|~(| dcache__GEN_55 )|~(| dcache__GEN_56 )|~(| dcache__GEN_58 )|~(| dcache__GEN_57 ); 
    wire[3:0] dcache_putpartial_mask = dcache_a_mask [3:0]; 
    wire dcache__atomics_legal_T_243 = dcache_s2_req_size !=2'h3; 
    wire[2:0] dcache__GEN_60 ={ dcache_s2_req_addr [30], dcache_s2_req_addr [27], dcache_s2_req_addr [16]}; 
    wire dcache_atomics_legal = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH ={ dcache_atomics_a_mask_sizeOH_shiftAmount ,1'h1}; 
    wire dcache_atomics_a_mask_size = dcache_atomics_a_mask_sizeOH [1]; 
    wire dcache_atomics_a_mask_eq_1 = dcache_atomics_a_mask_bit ; 
    wire dcache_atomics_a_mask_nbit =~ dcache_atomics_a_mask_bit ; 
    wire dcache_atomics_a_mask_eq = dcache_atomics_a_mask_nbit ; 
    wire dcache_atomics_a_mask_acc = dcache_s2_req_size [1]| dcache_atomics_a_mask_size & dcache_atomics_a_mask_eq ; 
    wire dcache_atomics_a_mask_acc_1 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size & dcache_atomics_a_mask_eq_1 ; 
    wire dcache_atomics_a_mask_size_1 = dcache_atomics_a_mask_sizeOH [0]; 
    wire dcache_atomics_a_mask_nbit_1 =~ dcache_atomics_a_mask_bit_1 ; 
    wire dcache_atomics_a_mask_eq_2 = dcache_atomics_a_mask_eq & dcache_atomics_a_mask_nbit_1 ; 
    wire dcache_atomics_a_mask_acc_2 = dcache_atomics_a_mask_acc | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_2 ; 
    wire dcache_atomics_a_mask_eq_3 = dcache_atomics_a_mask_eq & dcache_atomics_a_mask_bit_1 ; 
    wire dcache_atomics_a_mask_acc_3 = dcache_atomics_a_mask_acc | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_3 ; 
    wire dcache_atomics_a_mask_eq_4 = dcache_atomics_a_mask_eq_1 & dcache_atomics_a_mask_nbit_1 ; 
    wire dcache_atomics_a_mask_acc_4 = dcache_atomics_a_mask_acc_1 | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_4 ; 
    wire dcache_atomics_a_mask_eq_5 = dcache_atomics_a_mask_eq_1 & dcache_atomics_a_mask_bit_1 ; 
    wire dcache_atomics_a_mask_acc_5 = dcache_atomics_a_mask_acc_1 | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_5 ; 
    wire[1:0] dcache_atomics_a_mask_lo ={ dcache_atomics_a_mask_acc_3 , dcache_atomics_a_mask_acc_2 }; 
    wire[1:0] dcache_atomics_a_mask_hi ={ dcache_atomics_a_mask_acc_5 , dcache_atomics_a_mask_acc_4 }; 
    wire[3:0] dcache_atomics_a_mask ={ dcache_atomics_a_mask_hi , dcache_atomics_a_mask_lo }; 
    wire dcache_atomics_legal_1 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_1 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_1 ,1'h1}; 
    wire dcache_atomics_a_mask_size_2 = dcache_atomics_a_mask_sizeOH_1 [1]; 
    wire dcache_atomics_a_mask_eq_7 = dcache_atomics_a_mask_bit_2 ; 
    wire dcache_atomics_a_mask_nbit_2 =~ dcache_atomics_a_mask_bit_2 ; 
    wire dcache_atomics_a_mask_eq_6 = dcache_atomics_a_mask_nbit_2 ; 
    wire dcache_atomics_a_mask_acc_6 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_6 ; 
    wire dcache_atomics_a_mask_acc_7 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_7 ; 
    wire dcache_atomics_a_mask_size_3 = dcache_atomics_a_mask_sizeOH_1 [0]; 
    wire dcache_atomics_a_mask_nbit_3 =~ dcache_atomics_a_mask_bit_3 ; 
    wire dcache_atomics_a_mask_eq_8 = dcache_atomics_a_mask_eq_6 & dcache_atomics_a_mask_nbit_3 ; 
    wire dcache_atomics_a_mask_acc_8 = dcache_atomics_a_mask_acc_6 | dcache_atomics_a_mask_size_3 & dcache_atomics_a_mask_eq_8 ; 
    wire dcache_atomics_a_mask_eq_9 = dcache_atomics_a_mask_eq_6 & dcache_atomics_a_mask_bit_3 ; 
    wire dcache_atomics_a_mask_acc_9 = dcache_atomics_a_mask_acc_6 | dcache_atomics_a_mask_size_3 & dcache_atomics_a_mask_eq_9 ; 
    wire dcache_atomics_a_mask_eq_10 = dcache_atomics_a_mask_eq_7 & dcache_atomics_a_mask_nbit_3 ; 
    wire dcache_atomics_a_mask_acc_10 = dcache_atomics_a_mask_acc_7 | dcache_atomics_a_mask_size_3 & dcache_atomics_a_mask_eq_10 ; 
    wire dcache_atomics_a_mask_eq_11 = dcache_atomics_a_mask_eq_7 & dcache_atomics_a_mask_bit_3 ; 
    wire dcache_atomics_a_mask_acc_11 = dcache_atomics_a_mask_acc_7 | dcache_atomics_a_mask_size_3 & dcache_atomics_a_mask_eq_11 ; 
    wire[1:0] dcache_atomics_a_mask_lo_1 ={ dcache_atomics_a_mask_acc_9 , dcache_atomics_a_mask_acc_8 }; 
    wire[1:0] dcache_atomics_a_mask_hi_1 ={ dcache_atomics_a_mask_acc_11 , dcache_atomics_a_mask_acc_10 }; 
    wire[3:0] dcache_atomics_a_1_mask ={ dcache_atomics_a_mask_hi_1 , dcache_atomics_a_mask_lo_1 }; 
    wire dcache_atomics_legal_2 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_2 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_2 ,1'h1}; 
    wire dcache_atomics_a_mask_size_4 = dcache_atomics_a_mask_sizeOH_2 [1]; 
    wire dcache_atomics_a_mask_eq_13 = dcache_atomics_a_mask_bit_4 ; 
    wire dcache_atomics_a_mask_nbit_4 =~ dcache_atomics_a_mask_bit_4 ; 
    wire dcache_atomics_a_mask_eq_12 = dcache_atomics_a_mask_nbit_4 ; 
    wire dcache_atomics_a_mask_acc_12 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_4 & dcache_atomics_a_mask_eq_12 ; 
    wire dcache_atomics_a_mask_acc_13 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_4 & dcache_atomics_a_mask_eq_13 ; 
    wire dcache_atomics_a_mask_size_5 = dcache_atomics_a_mask_sizeOH_2 [0]; 
    wire dcache_atomics_a_mask_nbit_5 =~ dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_eq_14 = dcache_atomics_a_mask_eq_12 & dcache_atomics_a_mask_nbit_5 ; 
    wire dcache_atomics_a_mask_acc_14 = dcache_atomics_a_mask_acc_12 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_14 ; 
    wire dcache_atomics_a_mask_eq_15 = dcache_atomics_a_mask_eq_12 & dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_acc_15 = dcache_atomics_a_mask_acc_12 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_15 ; 
    wire dcache_atomics_a_mask_eq_16 = dcache_atomics_a_mask_eq_13 & dcache_atomics_a_mask_nbit_5 ; 
    wire dcache_atomics_a_mask_acc_16 = dcache_atomics_a_mask_acc_13 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_16 ; 
    wire dcache_atomics_a_mask_eq_17 = dcache_atomics_a_mask_eq_13 & dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_acc_17 = dcache_atomics_a_mask_acc_13 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_17 ; 
    wire[1:0] dcache_atomics_a_mask_lo_2 ={ dcache_atomics_a_mask_acc_15 , dcache_atomics_a_mask_acc_14 }; 
    wire[1:0] dcache_atomics_a_mask_hi_2 ={ dcache_atomics_a_mask_acc_17 , dcache_atomics_a_mask_acc_16 }; 
    wire[3:0] dcache_atomics_a_2_mask ={ dcache_atomics_a_mask_hi_2 , dcache_atomics_a_mask_lo_2 }; 
    wire dcache_atomics_legal_3 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_3 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_3 ,1'h1}; 
    wire dcache_atomics_a_mask_size_6 = dcache_atomics_a_mask_sizeOH_3 [1]; 
    wire dcache_atomics_a_mask_eq_19 = dcache_atomics_a_mask_bit_6 ; 
    wire dcache_atomics_a_mask_nbit_6 =~ dcache_atomics_a_mask_bit_6 ; 
    wire dcache_atomics_a_mask_eq_18 = dcache_atomics_a_mask_nbit_6 ; 
    wire dcache_atomics_a_mask_acc_18 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_6 & dcache_atomics_a_mask_eq_18 ; 
    wire dcache_atomics_a_mask_acc_19 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_6 & dcache_atomics_a_mask_eq_19 ; 
    wire dcache_atomics_a_mask_size_7 = dcache_atomics_a_mask_sizeOH_3 [0]; 
    wire dcache_atomics_a_mask_nbit_7 =~ dcache_atomics_a_mask_bit_7 ; 
    wire dcache_atomics_a_mask_eq_20 = dcache_atomics_a_mask_eq_18 & dcache_atomics_a_mask_nbit_7 ; 
    wire dcache_atomics_a_mask_acc_20 = dcache_atomics_a_mask_acc_18 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_20 ; 
    wire dcache_atomics_a_mask_eq_21 = dcache_atomics_a_mask_eq_18 & dcache_atomics_a_mask_bit_7 ; 
    wire dcache_atomics_a_mask_acc_21 = dcache_atomics_a_mask_acc_18 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_21 ; 
    wire dcache_atomics_a_mask_eq_22 = dcache_atomics_a_mask_eq_19 & dcache_atomics_a_mask_nbit_7 ; 
    wire dcache_atomics_a_mask_acc_22 = dcache_atomics_a_mask_acc_19 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_22 ; 
    wire dcache_atomics_a_mask_eq_23 = dcache_atomics_a_mask_eq_19 & dcache_atomics_a_mask_bit_7 ; 
    wire dcache_atomics_a_mask_acc_23 = dcache_atomics_a_mask_acc_19 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_23 ; 
    wire[1:0] dcache_atomics_a_mask_lo_3 ={ dcache_atomics_a_mask_acc_21 , dcache_atomics_a_mask_acc_20 }; 
    wire[1:0] dcache_atomics_a_mask_hi_3 ={ dcache_atomics_a_mask_acc_23 , dcache_atomics_a_mask_acc_22 }; 
    wire[3:0] dcache_atomics_a_3_mask ={ dcache_atomics_a_mask_hi_3 , dcache_atomics_a_mask_lo_3 }; 
    wire dcache_atomics_legal_4 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_4 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_4 ,1'h1}; 
    wire dcache_atomics_a_mask_size_8 = dcache_atomics_a_mask_sizeOH_4 [1]; 
    wire dcache_atomics_a_mask_eq_25 = dcache_atomics_a_mask_bit_8 ; 
    wire dcache_atomics_a_mask_nbit_8 =~ dcache_atomics_a_mask_bit_8 ; 
    wire dcache_atomics_a_mask_eq_24 = dcache_atomics_a_mask_nbit_8 ; 
    wire dcache_atomics_a_mask_acc_24 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_24 ; 
    wire dcache_atomics_a_mask_acc_25 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_25 ; 
    wire dcache_atomics_a_mask_size_9 = dcache_atomics_a_mask_sizeOH_4 [0]; 
    wire dcache_atomics_a_mask_nbit_9 =~ dcache_atomics_a_mask_bit_9 ; 
    wire dcache_atomics_a_mask_eq_26 = dcache_atomics_a_mask_eq_24 & dcache_atomics_a_mask_nbit_9 ; 
    wire dcache_atomics_a_mask_acc_26 = dcache_atomics_a_mask_acc_24 | dcache_atomics_a_mask_size_9 & dcache_atomics_a_mask_eq_26 ; 
    wire dcache_atomics_a_mask_eq_27 = dcache_atomics_a_mask_eq_24 & dcache_atomics_a_mask_bit_9 ; 
    wire dcache_atomics_a_mask_acc_27 = dcache_atomics_a_mask_acc_24 | dcache_atomics_a_mask_size_9 & dcache_atomics_a_mask_eq_27 ; 
    wire dcache_atomics_a_mask_eq_28 = dcache_atomics_a_mask_eq_25 & dcache_atomics_a_mask_nbit_9 ; 
    wire dcache_atomics_a_mask_acc_28 = dcache_atomics_a_mask_acc_25 | dcache_atomics_a_mask_size_9 & dcache_atomics_a_mask_eq_28 ; 
    wire dcache_atomics_a_mask_eq_29 = dcache_atomics_a_mask_eq_25 & dcache_atomics_a_mask_bit_9 ; 
    wire dcache_atomics_a_mask_acc_29 = dcache_atomics_a_mask_acc_25 | dcache_atomics_a_mask_size_9 & dcache_atomics_a_mask_eq_29 ; 
    wire[1:0] dcache_atomics_a_mask_lo_4 ={ dcache_atomics_a_mask_acc_27 , dcache_atomics_a_mask_acc_26 }; 
    wire[1:0] dcache_atomics_a_mask_hi_4 ={ dcache_atomics_a_mask_acc_29 , dcache_atomics_a_mask_acc_28 }; 
    wire[3:0] dcache_atomics_a_4_mask ={ dcache_atomics_a_mask_hi_4 , dcache_atomics_a_mask_lo_4 }; 
    wire dcache_atomics_legal_5 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_5 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_5 ,1'h1}; 
    wire dcache_atomics_a_mask_size_10 = dcache_atomics_a_mask_sizeOH_5 [1]; 
    wire dcache_atomics_a_mask_eq_31 = dcache_atomics_a_mask_bit_10 ; 
    wire dcache_atomics_a_mask_nbit_10 =~ dcache_atomics_a_mask_bit_10 ; 
    wire dcache_atomics_a_mask_eq_30 = dcache_atomics_a_mask_nbit_10 ; 
    wire dcache_atomics_a_mask_acc_30 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_10 & dcache_atomics_a_mask_eq_30 ; 
    wire dcache_atomics_a_mask_acc_31 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_10 & dcache_atomics_a_mask_eq_31 ; 
    wire dcache_atomics_a_mask_size_11 = dcache_atomics_a_mask_sizeOH_5 [0]; 
    wire dcache_atomics_a_mask_nbit_11 =~ dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_eq_32 = dcache_atomics_a_mask_eq_30 & dcache_atomics_a_mask_nbit_11 ; 
    wire dcache_atomics_a_mask_acc_32 = dcache_atomics_a_mask_acc_30 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_32 ; 
    wire dcache_atomics_a_mask_eq_33 = dcache_atomics_a_mask_eq_30 & dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_acc_33 = dcache_atomics_a_mask_acc_30 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_33 ; 
    wire dcache_atomics_a_mask_eq_34 = dcache_atomics_a_mask_eq_31 & dcache_atomics_a_mask_nbit_11 ; 
    wire dcache_atomics_a_mask_acc_34 = dcache_atomics_a_mask_acc_31 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_34 ; 
    wire dcache_atomics_a_mask_eq_35 = dcache_atomics_a_mask_eq_31 & dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_acc_35 = dcache_atomics_a_mask_acc_31 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_35 ; 
    wire[1:0] dcache_atomics_a_mask_lo_5 ={ dcache_atomics_a_mask_acc_33 , dcache_atomics_a_mask_acc_32 }; 
    wire[1:0] dcache_atomics_a_mask_hi_5 ={ dcache_atomics_a_mask_acc_35 , dcache_atomics_a_mask_acc_34 }; 
    wire[3:0] dcache_atomics_a_5_mask ={ dcache_atomics_a_mask_hi_5 , dcache_atomics_a_mask_lo_5 }; 
    wire dcache_atomics_legal_6 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_6 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_6 ,1'h1}; 
    wire dcache_atomics_a_mask_size_12 = dcache_atomics_a_mask_sizeOH_6 [1]; 
    wire dcache_atomics_a_mask_eq_37 = dcache_atomics_a_mask_bit_12 ; 
    wire dcache_atomics_a_mask_nbit_12 =~ dcache_atomics_a_mask_bit_12 ; 
    wire dcache_atomics_a_mask_eq_36 = dcache_atomics_a_mask_nbit_12 ; 
    wire dcache_atomics_a_mask_acc_36 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_12 & dcache_atomics_a_mask_eq_36 ; 
    wire dcache_atomics_a_mask_acc_37 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_12 & dcache_atomics_a_mask_eq_37 ; 
    wire dcache_atomics_a_mask_size_13 = dcache_atomics_a_mask_sizeOH_6 [0]; 
    wire dcache_atomics_a_mask_nbit_13 =~ dcache_atomics_a_mask_bit_13 ; 
    wire dcache_atomics_a_mask_eq_38 = dcache_atomics_a_mask_eq_36 & dcache_atomics_a_mask_nbit_13 ; 
    wire dcache_atomics_a_mask_acc_38 = dcache_atomics_a_mask_acc_36 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_38 ; 
    wire dcache_atomics_a_mask_eq_39 = dcache_atomics_a_mask_eq_36 & dcache_atomics_a_mask_bit_13 ; 
    wire dcache_atomics_a_mask_acc_39 = dcache_atomics_a_mask_acc_36 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_39 ; 
    wire dcache_atomics_a_mask_eq_40 = dcache_atomics_a_mask_eq_37 & dcache_atomics_a_mask_nbit_13 ; 
    wire dcache_atomics_a_mask_acc_40 = dcache_atomics_a_mask_acc_37 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_40 ; 
    wire dcache_atomics_a_mask_eq_41 = dcache_atomics_a_mask_eq_37 & dcache_atomics_a_mask_bit_13 ; 
    wire dcache_atomics_a_mask_acc_41 = dcache_atomics_a_mask_acc_37 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_41 ; 
    wire[1:0] dcache_atomics_a_mask_lo_6 ={ dcache_atomics_a_mask_acc_39 , dcache_atomics_a_mask_acc_38 }; 
    wire[1:0] dcache_atomics_a_mask_hi_6 ={ dcache_atomics_a_mask_acc_41 , dcache_atomics_a_mask_acc_40 }; 
    wire[3:0] dcache_atomics_a_6_mask ={ dcache_atomics_a_mask_hi_6 , dcache_atomics_a_mask_lo_6 }; 
    wire dcache_atomics_legal_7 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_7 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_7 ,1'h1}; 
    wire dcache_atomics_a_mask_size_14 = dcache_atomics_a_mask_sizeOH_7 [1]; 
    wire dcache_atomics_a_mask_eq_43 = dcache_atomics_a_mask_bit_14 ; 
    wire dcache_atomics_a_mask_nbit_14 =~ dcache_atomics_a_mask_bit_14 ; 
    wire dcache_atomics_a_mask_eq_42 = dcache_atomics_a_mask_nbit_14 ; 
    wire dcache_atomics_a_mask_acc_42 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_42 ; 
    wire dcache_atomics_a_mask_acc_43 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_43 ; 
    wire dcache_atomics_a_mask_size_15 = dcache_atomics_a_mask_sizeOH_7 [0]; 
    wire dcache_atomics_a_mask_nbit_15 =~ dcache_atomics_a_mask_bit_15 ; 
    wire dcache_atomics_a_mask_eq_44 = dcache_atomics_a_mask_eq_42 & dcache_atomics_a_mask_nbit_15 ; 
    wire dcache_atomics_a_mask_acc_44 = dcache_atomics_a_mask_acc_42 | dcache_atomics_a_mask_size_15 & dcache_atomics_a_mask_eq_44 ; 
    wire dcache_atomics_a_mask_eq_45 = dcache_atomics_a_mask_eq_42 & dcache_atomics_a_mask_bit_15 ; 
    wire dcache_atomics_a_mask_acc_45 = dcache_atomics_a_mask_acc_42 | dcache_atomics_a_mask_size_15 & dcache_atomics_a_mask_eq_45 ; 
    wire dcache_atomics_a_mask_eq_46 = dcache_atomics_a_mask_eq_43 & dcache_atomics_a_mask_nbit_15 ; 
    wire dcache_atomics_a_mask_acc_46 = dcache_atomics_a_mask_acc_43 | dcache_atomics_a_mask_size_15 & dcache_atomics_a_mask_eq_46 ; 
    wire dcache_atomics_a_mask_eq_47 = dcache_atomics_a_mask_eq_43 & dcache_atomics_a_mask_bit_15 ; 
    wire dcache_atomics_a_mask_acc_47 = dcache_atomics_a_mask_acc_43 | dcache_atomics_a_mask_size_15 & dcache_atomics_a_mask_eq_47 ; 
    wire[1:0] dcache_atomics_a_mask_lo_7 ={ dcache_atomics_a_mask_acc_45 , dcache_atomics_a_mask_acc_44 }; 
    wire[1:0] dcache_atomics_a_mask_hi_7 ={ dcache_atomics_a_mask_acc_47 , dcache_atomics_a_mask_acc_46 }; 
    wire[3:0] dcache_atomics_a_7_mask ={ dcache_atomics_a_mask_hi_7 , dcache_atomics_a_mask_lo_7 }; 
    wire dcache_atomics_legal_8 = dcache__atomics_legal_T_243 &(~(| dcache__GEN_60 )|~(| dcache__GEN_56 )); 
    wire[1:0] dcache_atomics_a_mask_sizeOH_8 ={ dcache_atomics_a_mask_sizeOH_shiftAmount_8 ,1'h1}; 
    wire dcache_atomics_a_mask_size_16 = dcache_atomics_a_mask_sizeOH_8 [1]; 
    wire dcache_atomics_a_mask_eq_49 = dcache_atomics_a_mask_bit_16 ; 
    wire dcache_atomics_a_mask_nbit_16 =~ dcache_atomics_a_mask_bit_16 ; 
    wire dcache_atomics_a_mask_eq_48 = dcache_atomics_a_mask_nbit_16 ; 
    wire dcache_atomics_a_mask_acc_48 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_16 & dcache_atomics_a_mask_eq_48 ; 
    wire dcache_atomics_a_mask_acc_49 = dcache_s2_req_size [1]| dcache_atomics_a_mask_size_16 & dcache_atomics_a_mask_eq_49 ; 
    wire dcache_atomics_a_mask_size_17 = dcache_atomics_a_mask_sizeOH_8 [0]; 
    wire dcache_atomics_a_mask_nbit_17 =~ dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_eq_50 = dcache_atomics_a_mask_eq_48 & dcache_atomics_a_mask_nbit_17 ; 
    wire dcache_atomics_a_mask_acc_50 = dcache_atomics_a_mask_acc_48 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_50 ; 
    wire dcache_atomics_a_mask_eq_51 = dcache_atomics_a_mask_eq_48 & dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_acc_51 = dcache_atomics_a_mask_acc_48 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_51 ; 
    wire dcache_atomics_a_mask_eq_52 = dcache_atomics_a_mask_eq_49 & dcache_atomics_a_mask_nbit_17 ; 
    wire dcache_atomics_a_mask_acc_52 = dcache_atomics_a_mask_acc_49 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_52 ; 
    wire dcache_atomics_a_mask_eq_53 = dcache_atomics_a_mask_eq_49 & dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_acc_53 = dcache_atomics_a_mask_acc_49 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_53 ; 
    wire[1:0] dcache_atomics_a_mask_lo_8 ={ dcache_atomics_a_mask_acc_51 , dcache_atomics_a_mask_acc_50 }; 
    wire[1:0] dcache_atomics_a_mask_hi_8 ={ dcache_atomics_a_mask_acc_53 , dcache_atomics_a_mask_acc_52 }; 
    wire[3:0] dcache_atomics_a_8_mask ={ dcache_atomics_a_mask_hi_8 , dcache_atomics_a_mask_lo_8 }; 
    wire dcache__atomics_T = dcache_s2_req_cmd ==5'h4; 
    wire dcache__atomics_T_2 = dcache_s2_req_cmd ==5'h9; 
    wire dcache__atomics_T_4 = dcache_s2_req_cmd ==5'hA; 
    wire dcache__atomics_T_6 = dcache_s2_req_cmd ==5'hB; 
    wire dcache__atomics_T_8 = dcache_s2_req_cmd ==5'h8; 
    wire dcache__atomics_T_10 = dcache_s2_req_cmd ==5'hC; 
    wire dcache__atomics_T_12 = dcache_s2_req_cmd ==5'hD; 
    wire dcache__atomics_T_14 = dcache_s2_req_cmd ==5'hE; 
    wire dcache__atomics_T_16 = dcache_s2_req_cmd ==5'hF; 
    wire[2:0] dcache_atomics_opcode = dcache__atomics_T_16 | dcache__atomics_T_14 | dcache__atomics_T_12 | dcache__atomics_T_10 | dcache__atomics_T_8  ? 3'h2: dcache__atomics_T_6 | dcache__atomics_T_4 | dcache__atomics_T_2 | dcache__atomics_T  ? 3'h3:3'h0; 
    wire[2:0] dcache_atomics_param = dcache__atomics_T_16  ? 3'h3: dcache__atomics_T_14  ? 3'h2: dcache__atomics_T_12  ? 3'h1: dcache__atomics_T_10  ? 3'h0: dcache__atomics_T_8  ? 3'h4: dcache__atomics_T_6  ? 3'h2: dcache__atomics_T_4  ? 3'h1: dcache__atomics_T_2 |~ dcache__atomics_T  ? 3'h0:3'h3; 
    wire[3:0] dcache_atomics_size = dcache__atomics_T_16  ?  dcache_atomics_a_8_size : dcache__atomics_T_14  ?  dcache_atomics_a_7_size : dcache__atomics_T_12  ?  dcache_atomics_a_6_size : dcache__atomics_T_10  ?  dcache_atomics_a_5_size : dcache__atomics_T_8  ?  dcache_atomics_a_4_size : dcache__atomics_T_6  ?  dcache_atomics_a_3_size : dcache__atomics_T_4  ?  dcache_atomics_a_2_size : dcache__atomics_T_2  ?  dcache_atomics_a_1_size : dcache__atomics_T  ?  dcache_atomics_a_size :4'h0; 
    wire[31:0] dcache_atomics_address = dcache__atomics_T_16  ?  dcache_atomics_a_8_address : dcache__atomics_T_14  ?  dcache_atomics_a_7_address : dcache__atomics_T_12  ?  dcache_atomics_a_6_address : dcache__atomics_T_10  ?  dcache_atomics_a_5_address : dcache__atomics_T_8  ?  dcache_atomics_a_4_address : dcache__atomics_T_6  ?  dcache_atomics_a_3_address : dcache__atomics_T_4  ?  dcache_atomics_a_2_address : dcache__atomics_T_2  ?  dcache_atomics_a_1_address : dcache__atomics_T  ?  dcache_atomics_a_address :32'h0; 
    wire[3:0] dcache_atomics_mask = dcache__atomics_T_16  ?  dcache_atomics_a_8_mask : dcache__atomics_T_14  ?  dcache_atomics_a_7_mask : dcache__atomics_T_12  ?  dcache_atomics_a_6_mask : dcache__atomics_T_10  ?  dcache_atomics_a_5_mask : dcache__atomics_T_8  ?  dcache_atomics_a_4_mask : dcache__atomics_T_6  ?  dcache_atomics_a_3_mask : dcache__atomics_T_4  ?  dcache_atomics_a_2_mask : dcache__atomics_T_2  ?  dcache_atomics_a_1_mask : dcache__atomics_T  ?  dcache_atomics_a_mask :4'h0; 
    wire[31:0] dcache_atomics_data = dcache__atomics_T_16  ?  dcache_atomics_a_8_data : dcache__atomics_T_14  ?  dcache_atomics_a_7_data : dcache__atomics_T_12  ?  dcache_atomics_a_6_data : dcache__atomics_T_10  ?  dcache_atomics_a_5_data : dcache__atomics_T_8  ?  dcache_atomics_a_4_data : dcache__atomics_T_6  ?  dcache_atomics_a_3_data : dcache__atomics_T_4  ?  dcache_atomics_a_2_data : dcache__atomics_T_2  ?  dcache_atomics_a_1_data : dcache__atomics_T  ?  dcache_atomics_a_data :32'h0; 
  assign  dcache_tl_out_a_valid = dcache_s2_valid_uncached_pending | dcache_s2_valid_cached_miss &~ dcache_s2_victim_dirty ; 
  assign  dcache_tl_out_a_bits_opcode = dcache_s2_uncached  ? ( dcache_s2_write  ? ( dcache__metaArb_io_in_3_bits_data_c_cat_T_24  ? 3'h1: dcache_s2_read  ?  dcache_atomics_opcode :3'h0):3'h4):3'h0; 
    wire dcache__GEN_61 =~ dcache_s2_uncached |~ dcache_s2_write ; 
  assign  dcache_tl_out_a_bits_param = dcache__GEN_61 | dcache__metaArb_io_in_3_bits_data_c_cat_T_24 |~ dcache_s2_read  ? 3'h0: dcache_atomics_param ; 
  assign  dcache_tl_out_a_bits_size = dcache_s2_uncached  ? ( dcache_s2_write  ? ( dcache__metaArb_io_in_3_bits_data_c_cat_T_24  ?  dcache_putpartial_size : dcache_s2_read  ?  dcache_atomics_size : dcache_put_size ): dcache_get_size ):4'h0; 
  assign  dcache_tl_out_a_bits_address = dcache_s2_uncached  ? ( dcache_s2_write  ? ( dcache__metaArb_io_in_3_bits_data_c_cat_T_24  ?  dcache_putpartial_address : dcache_s2_read  ?  dcache_atomics_address : dcache_put_address ): dcache_get_address ):32'h0; 
  assign  dcache_tl_out_a_bits_mask = dcache_s2_uncached  ? ( dcache_s2_write  ? ( dcache__metaArb_io_in_3_bits_data_c_cat_T_24  ?  dcache_putpartial_mask : dcache_s2_read  ?  dcache_atomics_mask : dcache_put_mask ): dcache_get_mask ):4'h0; 
  assign  dcache_tl_out_a_bits_data = dcache__GEN_61  ? 32'h0: dcache__metaArb_io_in_3_bits_data_c_cat_T_24  ?  dcache_putpartial_data : dcache_s2_read  ?  dcache_atomics_data : dcache_put_data ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_privileged =(& dcache_s2_req_dprv )| dcache_s2_pma_cacheable ; 
    wire dcache__io_cpu_perf_acquire_T = dcache_tl_out_a_ready & dcache_tl_out_a_valid ; 
    wire dcache_nodeOut_d_ready ; 
    wire dcache__io_errors_bus_valid_T = dcache_nodeOut_d_ready & dcache_nodeOut_d_valid ; 
    wire[26:0] dcache__beats1_decode_T_1 =27'hFFF<< dcache_nodeOut_d_bits_size ; 
    wire[9:0] dcache_beats1_decode =~( dcache__beats1_decode_T_1 [11:2]); 
    wire dcache_beats1_opdata = dcache_nodeOut_d_bits_opcode [0]; 
    wire[9:0] dcache_beats1 = dcache_beats1_opdata  ?  dcache_beats1_decode :10'h0; reg[9:0] dcache_counter ; 
    wire[9:0] dcache_counter1 = dcache_counter -10'h1; 
    wire dcache_d_first = dcache_counter ==10'h0; 
    wire dcache_d_last = dcache_counter ==10'h1| dcache_beats1 ==10'h0; 
    wire dcache_d_done = dcache_d_last & dcache__io_errors_bus_valid_T ; 
    wire[9:0] dcache_count = dcache_beats1 &~ dcache_counter1 ; 
    wire[11:0] dcache_d_address_inc ={ dcache_count ,2'h0}; 
    wire[1:0] dcache_d_opc = dcache_nodeOut_d_bits_opcode [1:0]; 
    wire[1:0] dcache_data_plaInput = dcache_d_opc ; 
    wire[1:0] dcache_data_invInputs =~ dcache_data_plaInput ; 
    wire dcache_data_invMatrixOutputs ; 
    wire dcache_grantIsUncachedData = dcache_data_plaOutput ; 
    wire dcache_data_andMatrixInput_0 = dcache_data_plaInput [0]; 
    wire dcache_data_andMatrixInput_1 = dcache_data_invInputs [1]; 
    wire dcache_data_orMatrixOutputs =&{ dcache_data_andMatrixInput_0 , dcache_data_andMatrixInput_1 }; 
  assign  dcache_data_invMatrixOutputs = dcache_data_orMatrixOutputs ; 
  assign  dcache_data_plaOutput = dcache_data_invMatrixOutputs ; 
  assign  dcache_tl_d_data_encoded ={ dcache_tl_d_data_encoded_hi_1 , dcache_tl_d_data_encoded_lo_1 }; 
    reg dcache_grantInProgress ; 
    wire dcache_block_probe_for_ordering = dcache_grantInProgress ; reg[2:0] dcache_blockProbeAfterGrantCount ; 
    wire dcache__GEN_62 = dcache__io_errors_bus_valid_T & dcache_grantIsCached ; 
    wire dcache_replace = dcache__GEN_62 & dcache_d_last ; 
    wire dcache__GEN_63 =~ dcache__io_errors_bus_valid_T | dcache_grantIsCached |~ dcache_grantIsUncachedData ; 
    wire[1:0] dcache_s1_data_way = dcache__GEN_63  ? 2'h1:2'h2; 
    wire[31:0] dcache_s2_req_addr_dontCareBits ={ dcache_s1_paddr [31:2],2'h0}; 
  assign  dcache_metaArb_io_in_3_valid = dcache_grantIsCached & dcache_d_done &~ dcache_nodeOut_d_bits_denied ; 
    wire[1:0] dcache_metaArb_io_in_3_bits_data_c ={ dcache__metaArb_io_in_3_bits_data_c_cat_T_23 | dcache__metaArb_io_in_3_bits_data_c_cat_T_24 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 | dcache__metaArb_io_in_3_bits_data_c_cat_T_28 | dcache__metaArb_io_in_3_bits_data_c_cat_T_29 | dcache__metaArb_io_in_3_bits_data_c_cat_T_30 | dcache__metaArb_io_in_3_bits_data_c_cat_T_31 | dcache__metaArb_io_in_3_bits_data_c_cat_T_35 | dcache__metaArb_io_in_3_bits_data_c_cat_T_36 | dcache__metaArb_io_in_3_bits_data_c_cat_T_37 | dcache__metaArb_io_in_3_bits_data_c_cat_T_38 | dcache__metaArb_io_in_3_bits_data_c_cat_T_39 , dcache__metaArb_io_in_3_bits_data_c_cat_T_23 | dcache__metaArb_io_in_3_bits_data_c_cat_T_24 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 | dcache__metaArb_io_in_3_bits_data_c_cat_T_28 | dcache__metaArb_io_in_3_bits_data_c_cat_T_29 | dcache__metaArb_io_in_3_bits_data_c_cat_T_30 | dcache__metaArb_io_in_3_bits_data_c_cat_T_31 | dcache__metaArb_io_in_3_bits_data_c_cat_T_35 | dcache__metaArb_io_in_3_bits_data_c_cat_T_36 | dcache__metaArb_io_in_3_bits_data_c_cat_T_37 | dcache__metaArb_io_in_3_bits_data_c_cat_T_38 | dcache__metaArb_io_in_3_bits_data_c_cat_T_39 | dcache__metaArb_io_in_3_bits_data_c_cat_T_46 | dcache__metaArb_io_in_3_bits_data_c_cat_T_48 }; 
    wire[3:0] dcache__metaArb_io_in_3_bits_data_T_1 ={ dcache_metaArb_io_in_3_bits_data_c , dcache_nodeOut_d_bits_param }; 
    wire[1:0] dcache_metaArb_io_in_3_bits_data_meta_state = dcache__metaArb_io_in_3_bits_data_T_1 ==4'hC ? 2'h3: dcache__metaArb_io_in_3_bits_data_T_1 ==4'h4| dcache__metaArb_io_in_3_bits_data_T_1 ==4'h0 ? 2'h2:{1'h0, dcache__metaArb_io_in_3_bits_data_T_1 ==4'h1}; 
    wire[1:0] dcache_metaArb_io_in_3_bits_data_meta_1_coh_state = dcache_metaArb_io_in_3_bits_data_meta_state ; 
    reg dcache_blockUncachedGrant ; 
    wire dcache__GEN_64 = dcache_grantIsUncachedData &( dcache_blockUncachedGrant | dcache_s1_valid ); 
  assign  dcache_nodeOut_d_ready =~( dcache__GEN_64 | dcache_grantIsRefill &~ dcache_dataArb_grant_1 )&(~ dcache_grantIsCached |~ dcache_d_first ); 
    wire dcache__io_cpu_req_ready_output = dcache__GEN_64  ? ~( dcache_nodeOut_d_valid | dcache__GEN_47 )& dcache__io_cpu_req_ready_T_4 :~ dcache__GEN_47 & dcache__io_cpu_req_ready_T_4 ; 
    wire dcache__GEN_65 = dcache__GEN_64 & dcache_nodeOut_d_valid ; 
  assign  dcache_dataArb_io_in_1_valid = dcache__GEN_65 | dcache_nodeOut_d_valid & dcache_grantIsRefill ; 
  assign  dcache__GEN =~ dcache__GEN_65 ; 
    wire dcache_block_probe_for_core_progress =(| dcache_blockProbeAfterGrantCount )| dcache_lrscValid ; 
    wire[3:0] dcache_tl_out_c_bits_size ; 
    wire[26:0] dcache__GEN_66 ={23'h0, dcache_tl_out_c_bits_size }; 
    wire[26:0] dcache__beats1_decode_T_5 =27'hFFF<< dcache__GEN_66 ; 
    wire[9:0] dcache_beats1_decode_1 =~( dcache__beats1_decode_T_5 [11:2]); 
    reg dcache_s2_release_data_valid ; 
    wire dcache_tl_out_c_valid = dcache_s2_release_data_valid ; 
    wire dcache_releaseRejected = dcache_s2_release_data_valid ; 
    wire[10:0] dcache_releaseDataBeat ={9'h0, dcache_releaseRejected  ? 2'h0:{1'h0, dcache_s2_release_data_valid }}; 
  assign  dcache_tl_out_c_bits_size = dcache_nackResponseMessage_size ; 
    wire dcache_tl_out_c_bits_source = dcache_nackResponseMessage_source ; 
    wire[31:0] dcache_tl_out_c_bits_address = dcache_nackResponseMessage_address ; 
    wire[1:0] dcache_metaArb_io_in_4_bits_data_meta_coh_state = dcache_newCoh_state ; 
    wire[17:0] dcache_metaArb_io_in_4_bits_data_meta_tag = dcache_tl_out_c_bits_address [31:14]; 
    wire dcache_s1_xcpt_valid = dcache_s1_valid &~ dcache_io_cpu_s1_kill & dcache_s1_cmd_uses_tlb &~ dcache_s1_req_no_xcpt &~ dcache_s1_nack ; 
    reg dcache_io_cpu_s2_xcpt_REG ; 
  assign  dcache__io_cpu_s2_xcpt_pf_ld_output = dcache_io_cpu_s2_xcpt_REG & dcache_s2_tlb_xcpt_pf_ld ; 
  assign  dcache__io_cpu_s2_xcpt_pf_st_output = dcache_io_cpu_s2_xcpt_REG & dcache_s2_tlb_xcpt_pf_st ; 
  assign  dcache__io_cpu_s2_xcpt_ae_ld_output = dcache_io_cpu_s2_xcpt_REG & dcache_s2_tlb_xcpt_ae_ld ; 
  assign  dcache__io_cpu_s2_xcpt_ae_st_output = dcache_io_cpu_s2_xcpt_REG & dcache_s2_tlb_xcpt_ae_st ; 
  assign  dcache__io_cpu_s2_xcpt_ma_ld_output = dcache_io_cpu_s2_xcpt_REG & dcache_s2_tlb_xcpt_ma_ld ; 
  assign  dcache__io_cpu_s2_xcpt_ma_st_output = dcache_io_cpu_s2_xcpt_REG & dcache_s2_tlb_xcpt_ma_st ; reg[31:0] dcache_s2_uncached_data_word ; 
    reg dcache_doUncachedResp ; 
  assign  dcache__io_cpu_replay_next_output = dcache__io_errors_bus_valid_T & dcache_grantIsUncachedData ; 
  always @( posedge  dcache_clock )
         begin 
             if (~ dcache_reset &~(~( dcache__pstore_drain_opportunistic_T | dcache__pstore_drain_opportunistic_T_1 | dcache__pstore_drain_opportunistic_T_2 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 |( dcache__pstore_drain_opportunistic_T_25 | dcache__pstore_drain_opportunistic_T_50 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 )& dcache__pstore_drain_opportunistic_T_50 )| dcache_dataArb_io_in_3_valid_res ))
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
                     if (1)$fatal;
                 end 
             if (~ dcache_reset &~(~( dcache_s1_valid_masked & dcache__io_cpu_perf_canAcceptLoadThenLoad_T_51 )|(&( dcache_s1_mask_xwr |~ dcache_io_cpu_s1_data_mask ))))
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:306 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n");
                     if (1)$fatal;
                 end 
             if (~ dcache_reset &~(~( dcache__pstore_drain_opportunistic_T | dcache__pstore_drain_opportunistic_T_1 | dcache__pstore_drain_opportunistic_T_2 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 |( dcache__pstore_drain_opportunistic_T_25 | dcache__pstore_drain_opportunistic_T_50 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 )& dcache__pstore_drain_opportunistic_T_50 )| dcache_pstore_drain_opportunistic_res ))
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
                     if (1)$fatal;
                 end 
             if (~ dcache_reset &~( dcache_pstore1_rmw |( dcache__dataArb_io_in_0_valid_T_2 | dcache_pstore1_held )== dcache_pstore1_valid ))
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:487 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n");
                     if (1)$fatal;
                 end 
             if (~ dcache_reset &~(~ dcache_nodeOut_d_valid | dcache_nodeOut_d_bits_opcode ==3'h1| dcache_nodeOut_d_bits_opcode ==3'h0| dcache_nodeOut_d_bits_opcode ==3'h2))
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:631 assert(!tl_out.d.valid || whole_opc.isOneOf(uncachedGrantOpcodes))\n");
                     if (1)$fatal;
                 end 
             if ( dcache__GEN_62 &~ dcache_reset &~ dcache_cached_grant_wait )
                 begin 
                     if (1)$error("Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:654 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n");
                     if (1)$fatal;
                 end 
             if ( dcache__io_errors_bus_valid_T &~ dcache_grantIsCached & dcache_d_last &~ dcache_reset &~ dcache_uncachedInFlight_0 )
                 begin 
                     if (1)$error("Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:664 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n");
                     if (1)$fatal;
                 end 
             if (~ dcache_reset & dcache__io_errors_bus_valid_T & dcache_d_first & dcache_grantIsCached )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:693 assert(tl_out.e.fire === (tl_out.d.fire && d_first && grantIsCached))\n");
                     if (1)$fatal;
                 end 
             if (~ dcache_reset & dcache_s2_valid_masked &( dcache__metaArb_io_in_3_bits_data_c_cat_T_48 | dcache__metaArb_io_in_3_bits_data_c_cat_T_26 ))
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:912 assert(!(s2_valid_masked && s2_req.cmd.isOneOf(M_XLR, M_XSC)))\n");
                     if (1)$fatal;
                 end 
             if ( dcache_doUncachedResp &~ dcache_reset & dcache_s2_valid_hit )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:928 assert(!s2_valid_hit)\n");
                     if (1)$fatal;
                 end 
         end
    wire[31:0] dcache_s2_data_word_possibly_uncached = dcache_s2_data_word ; 
    wire[15:0] dcache_io_cpu_resp_bits_data_shifted = dcache_s2_req_addr [1] ?  dcache_s2_data_word_possibly_uncached [31:16]: dcache_s2_data_word_possibly_uncached [15:0]; 
    wire[15:0] dcache_io_cpu_resp_bits_data_zeroed = dcache_io_cpu_resp_bits_data_shifted ; 
    wire[7:0] dcache_io_cpu_resp_bits_data_shifted_1 = dcache_s2_req_addr [0] ?  dcache_io_cpu_resp_bits_data_zeroed [15:8]: dcache_io_cpu_resp_bits_data_zeroed [7:0]; 
    wire[7:0] dcache_io_cpu_resp_bits_data_zeroed_1 = dcache_io_cpu_resp_bits_data_shifted_1 ; 
    wire[15:0] dcache_pstore1_storegen_data_mask_lo ={{8{ dcache_pstore1_mask [1]}},{8{ dcache_pstore1_mask [0]}}}; 
    wire[15:0] dcache_pstore1_storegen_data_mask_hi ={{8{ dcache_pstore1_mask [3]}},{8{ dcache_pstore1_mask [2]}}}; 
    wire[31:0] dcache_pstore1_storegen_data_mask ={ dcache_pstore1_storegen_data_mask_hi , dcache_pstore1_storegen_data_mask_lo }; 
    wire[31:0] dcache_pstore1_storegen_data = dcache__amoalus_0_io_out_unmasked & dcache_pstore1_storegen_data_mask | dcache_s2_data_word_corrected &~ dcache_pstore1_storegen_data_mask ; 
    wire[26:0] dcache__io_cpu_perf_acquire_beats1_decode_T_1 =27'hFFF<< dcache_tl_out_a_bits_size ; 
    wire[9:0] dcache_io_cpu_perf_acquire_beats1_decode =~( dcache__io_cpu_perf_acquire_beats1_decode_T_1 [11:2]); 
    wire dcache_io_cpu_perf_acquire_beats1_opdata =~( dcache_tl_out_a_bits_opcode [2]); 
    wire[9:0] dcache_io_cpu_perf_acquire_beats1 = dcache_io_cpu_perf_acquire_beats1_opdata  ?  dcache_io_cpu_perf_acquire_beats1_decode :10'h0; reg[9:0] dcache_io_cpu_perf_acquire_counter ; 
    wire[9:0] dcache_io_cpu_perf_acquire_counter1 = dcache_io_cpu_perf_acquire_counter -10'h1; 
    wire dcache_io_cpu_perf_acquire_first = dcache_io_cpu_perf_acquire_counter ==10'h0; 
    wire dcache_io_cpu_perf_acquire_last = dcache_io_cpu_perf_acquire_counter ==10'h1| dcache_io_cpu_perf_acquire_beats1 ==10'h0; 
    wire dcache_io_cpu_perf_acquire_done = dcache_io_cpu_perf_acquire_last & dcache__io_cpu_perf_acquire_T ; 
    wire[9:0] dcache_io_cpu_perf_acquire_count = dcache_io_cpu_perf_acquire_beats1 &~ dcache_io_cpu_perf_acquire_counter1 ; 
    wire[26:0] dcache__io_cpu_perf_release_beats1_decode_T_1 =27'hFFF<< dcache__GEN_66 ; 
    wire[9:0] dcache_io_cpu_perf_release_beats1_decode =~( dcache__io_cpu_perf_release_beats1_decode_T_1 [11:2]); reg[3:0] dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count ; 
    wire dcache_io_cpu_perf_blocked_near_end_of_refill = dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count >4'hD; 
    wire dcache__GEN_67 = dcache__io_errors_bus_valid_T & dcache_grantIsCached & dcache_d_last ; 
    wire dcache_tlb_io_resp_ma_ld = dcache_tlb_misaligned & dcache_tlb_cmd_read ; 
    wire dcache_tlb_io_resp_ma_st = dcache_tlb_misaligned & dcache_tlb_cmd_write ; 
    wire[31:0] dcache_tlb_io_resp_paddr ={ dcache_tlb_ppn , dcache_tlb_io_resp_gpa_offset }; 
    wire[31:0] dcache_tlb_io_resp_gpa ={ dcache_tlb_io_resp_gpa_page [19:0], dcache_tlb_io_resp_gpa_offset }; 
    wire[1:0] dcache__s2_data_T_1 = dcache_s2_data_s1_word_en  ?  dcache_s1_data_way :2'h0; 
    wire dcache__GEN_68 = dcache__io_cpu_perf_acquire_T & dcache_s2_uncached ; 
  always @( posedge  dcache_clock )
         begin 
             if ( dcache_reset )
                 begin  
                     dcache_s1_valid  <=1'h0; 
                     dcache_cached_grant_wait  <=1'h0; 
                     dcache_uncachedInFlight_0  <=1'h0; 
                     dcache_s2_valid  <=1'h0; 
                     dcache_lrscCount  <=7'h0; 
                     dcache_pstore2_valid  <=1'h0; 
                     dcache_pstore1_held  <=1'h0; 
                     dcache_counter  <=10'h0; 
                     dcache_grantInProgress  <=1'h0; 
                     dcache_blockProbeAfterGrantCount  <=3'h0; 
                     dcache_io_cpu_perf_acquire_counter  <=10'h0; 
                     dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count  <=4'h0;
                 end 
              else 
                 begin  
                     dcache_s1_valid  <= dcache__io_cpu_req_ready_output & dcache_io_cpu_req_valid ; 
                     dcache_cached_grant_wait  <=~ dcache__GEN_67 &( dcache__io_cpu_perf_acquire_T &~ dcache_s2_uncached | dcache_cached_grant_wait ); 
                     dcache_uncachedInFlight_0  <=(~ dcache__io_errors_bus_valid_T | dcache_grantIsCached |~ dcache_d_last )&( dcache__GEN_68 | dcache_uncachedInFlight_0 ); 
                     dcache_s2_valid  <= dcache_s1_valid_masked &~ dcache_s1_sfence ;
                     if ( dcache_s2_valid_not_killed & dcache_lrscValid ) 
                         dcache_lrscCount  <=7'h3;
                      else 
                         if (| dcache_lrscCount ) 
                             dcache_lrscCount  <= dcache_lrscCount -7'h1;
                          else 
                             if ( dcache_s2_valid_cached_miss ) 
                                 dcache_lrscCount  <= dcache_s2_hit  ? 7'h4F:7'h0; 
                     dcache_pstore2_valid  <= dcache_pstore2_valid &~ dcache_pstore_drain | dcache_advance_pstore1 ; 
                     dcache_pstore1_held  <=( dcache__pstore1_held_T | dcache_pstore1_held )& dcache_pstore2_valid &~ dcache_pstore_drain ;
                     if ( dcache__io_errors_bus_valid_T )
                         begin 
                             if ( dcache_d_first ) 
                                 dcache_counter  <= dcache_beats1 ;
                              else  
                                 dcache_counter  <= dcache_counter1 ;
                         end 
                     if ( dcache__GEN_62 ) 
                         dcache_grantInProgress  <=~ dcache_d_last ;
                     if ( dcache__GEN_67 ) 
                         dcache_blockProbeAfterGrantCount  <=3'h7;
                      else 
                         if (| dcache_blockProbeAfterGrantCount ) 
                             dcache_blockProbeAfterGrantCount  <= dcache_blockProbeAfterGrantCount -3'h1;
                     if ( dcache__io_cpu_perf_acquire_T )
                         begin 
                             if ( dcache_io_cpu_perf_acquire_first ) 
                                 dcache_io_cpu_perf_acquire_counter  <= dcache_io_cpu_perf_acquire_beats1 ;
                              else  
                                 dcache_io_cpu_perf_acquire_counter  <= dcache_io_cpu_perf_acquire_counter1 ;
                         end 
                     if ( dcache__io_errors_bus_valid_T & dcache_grantIsRefill ) 
                         dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count  <= dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count +4'h1;
                 end 
             if ( dcache_s0_clk_en )
                 begin  
                     dcache_s1_req_addr  <= dcache_s0_req_addr ; 
                     dcache_s1_req_tag  <= dcache_s0_req_tag ; 
                     dcache_s1_req_cmd  <= dcache_s0_req_cmd ; 
                     dcache_s1_req_size  <= dcache_s0_req_size ; 
                     dcache_s1_req_signed  <= dcache_s0_req_signed ; 
                     dcache_s1_req_dprv  <= dcache_s0_req_dprv ; 
                     dcache_s1_req_dv  <= dcache_s0_req_dv ; 
                     dcache_s1_req_phys  <= dcache_s0_req_phys ; 
                     dcache_s1_req_no_xcpt  <= dcache_s0_req_no_xcpt ; 
                     dcache_s1_tlb_req_vaddr  <= dcache_s0_tlb_req_vaddr ; 
                     dcache_s1_tlb_req_passthrough  <= dcache_s0_tlb_req_passthrough ; 
                     dcache_s1_tlb_req_size  <= dcache_s0_tlb_req_size ; 
                     dcache_s1_tlb_req_cmd  <= dcache_s0_tlb_req_cmd ; 
                     dcache_s1_tlb_req_prv  <= dcache_s0_tlb_req_prv ; 
                     dcache_s1_tlb_req_v  <= dcache_s0_tlb_req_v ; 
                     dcache_s1_did_read  <= dcache_dataArb_grant_3 & dcache_io_cpu_req_valid &( dcache__pstore_drain_opportunistic_T | dcache__pstore_drain_opportunistic_T_1 | dcache__pstore_drain_opportunistic_T_2 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 |( dcache__pstore_drain_opportunistic_T_25 | dcache__pstore_drain_opportunistic_T_50 | dcache__pstore_drain_opportunistic_T_28 | dcache__pstore_drain_opportunistic_T_30 | dcache__pstore_drain_opportunistic_T_31 | dcache__pstore_drain_opportunistic_T_32 | dcache__pstore_drain_opportunistic_T_33 | dcache__pstore_drain_opportunistic_T_37 | dcache__pstore_drain_opportunistic_T_38 | dcache__pstore_drain_opportunistic_T_39 | dcache__pstore_drain_opportunistic_T_40 | dcache__pstore_drain_opportunistic_T_41 )& dcache__pstore_drain_opportunistic_T_50 );
                 end  
             dcache_s1_flush_valid  <=1'h0;
             if (~ dcache__io_cpu_perf_acquire_T | dcache_s2_uncached )
                 begin 
                 end 
              else  
                 dcache_refill_way  <= dcache_s2_victim_or_hit_way ;
             if ( dcache__GEN_68 )
                 begin  
                     dcache_uncachedReqs_0_addr  <= dcache_s2_req_addr ; 
                     dcache_uncachedReqs_0_tag  <= dcache_s2_req_tag ; 
                     dcache_uncachedReqs_0_cmd  <= dcache_s2_write  ? { dcache__metaArb_io_in_3_bits_data_c_cat_T_24 ,4'h1}:5'h0; 
                     dcache_uncachedReqs_0_size  <= dcache_s2_req_size ; 
                     dcache_uncachedReqs_0_signed  <= dcache_s2_req_signed ; 
                     dcache_uncachedReqs_0_dprv  <= dcache_s2_req_dprv ; 
                     dcache_uncachedReqs_0_dv  <= dcache_s2_req_dv ; 
                     dcache_uncachedReqs_0_phys  <= dcache_s2_req_phys ; 
                     dcache_uncachedReqs_0_no_alloc  <= dcache_s2_req_no_alloc ; 
                     dcache_uncachedReqs_0_no_xcpt  <= dcache_s2_req_no_xcpt ; 
                     dcache_uncachedReqs_0_data  <= dcache_s2_req_data ; 
                     dcache_uncachedReqs_0_mask  <= dcache_s2_req_mask ;
                 end  
             dcache_s2_not_nacked_in_s1  <=~ dcache_s1_nack ;
             if ( dcache__GEN_63 )
                 begin 
                     if ( dcache_s1_meta_clk_en )
                         begin  
                             dcache_s2_req_addr  <= dcache_s1_paddr ; 
                             dcache_s2_req_tag  <= dcache_s1_req_tag ; 
                             dcache_s2_req_cmd  <= dcache_s1_req_cmd ; 
                             dcache_s2_req_size  <= dcache_s1_req_size ; 
                             dcache_s2_req_signed  <= dcache_s1_req_signed ;
                         end 
                 end 
              else 
                 begin  
                     dcache_s2_req_addr  <={ dcache_s2_req_addr_dontCareBits [31:2], dcache_s2_req_addr_dontCareBits [1:0]| dcache_uncachedResp_addr [1:0]}; 
                     dcache_s2_req_tag  <= dcache_uncachedResp_tag ; 
                     dcache_s2_req_cmd  <=5'h0; 
                     dcache_s2_req_size  <= dcache_uncachedResp_size ; 
                     dcache_s2_req_signed  <= dcache_uncachedResp_signed ;
                 end 
             if ( dcache_s1_meta_clk_en )
                 begin  
                     dcache_s2_req_dprv  <= dcache_s1_req_dprv ; 
                     dcache_s2_req_dv  <= dcache_s1_req_dv ; 
                     dcache_s2_req_phys  <= dcache_s1_req_phys ; 
                     dcache_s2_req_no_xcpt  <= dcache_s1_req_no_xcpt ; 
                     dcache_s2_req_data  <=32'h0; 
                     dcache_s2_req_mask  <=4'h0; 
                     dcache_s2_tlb_xcpt_paddr  <= dcache_tlb_io_resp_paddr ; 
                     dcache_s2_tlb_xcpt_gpa  <= dcache_tlb_io_resp_gpa ; 
                     dcache_s2_tlb_xcpt_pf_ld  <= dcache_tlb_pf_ld_array [6]; 
                     dcache_s2_tlb_xcpt_pf_st  <= dcache_tlb_pf_st_array [6]; 
                     dcache_s2_tlb_xcpt_pf_inst  <= dcache_tlb_pf_inst_array [6]; 
                     dcache_s2_tlb_xcpt_ae_ld  <= dcache_tlb_ae_ld_array [6]; 
                     dcache_s2_tlb_xcpt_ae_st  <= dcache_tlb_ae_st_array [6]; 
                     dcache_s2_tlb_xcpt_ae_inst  <=~( dcache_tlb_px_array [6]); 
                     dcache_s2_tlb_xcpt_ma_ld  <= dcache_tlb_io_resp_ma_ld ; 
                     dcache_s2_tlb_xcpt_ma_st  <= dcache_tlb_io_resp_ma_st ; 
                     dcache_s2_tlb_xcpt_cacheable  <= dcache_tlb_c_array [6]; 
                     dcache_s2_tlb_xcpt_must_alloc  <= dcache_tlb_must_alloc_array [6]; 
                     dcache_s2_tlb_xcpt_prefetchable  <= dcache_tlb_prefetchable_array [6]; 
                     dcache_s2_pma_paddr  <= dcache_tlb_io_resp_paddr ; 
                     dcache_s2_pma_gpa  <= dcache_tlb_io_resp_gpa ; 
                     dcache_s2_pma_pf_ld  <= dcache_tlb_pf_ld_array [6]; 
                     dcache_s2_pma_pf_st  <= dcache_tlb_pf_st_array [6]; 
                     dcache_s2_pma_pf_inst  <= dcache_tlb_pf_inst_array [6]; 
                     dcache_s2_pma_ae_ld  <= dcache_tlb_ae_ld_array [6]; 
                     dcache_s2_pma_ae_st  <= dcache_tlb_ae_st_array [6]; 
                     dcache_s2_pma_ae_inst  <=~( dcache_tlb_px_array [6]); 
                     dcache_s2_pma_ma_ld  <= dcache_tlb_io_resp_ma_ld ; 
                     dcache_s2_pma_ma_st  <= dcache_tlb_io_resp_ma_st ; 
                     dcache_s2_pma_cacheable  <= dcache_tlb_c_array [6]; 
                     dcache_s2_pma_must_alloc  <= dcache_tlb_must_alloc_array [6]; 
                     dcache_s2_pma_prefetchable  <= dcache_tlb_prefetchable_array [6]; 
                     dcache_s2_vaddr_r  <= dcache_s1_vaddr ; 
                     dcache_s2_hit_state_state  <= dcache_s1_hit_state_state ;
                 end  
             dcache_s2_req_no_alloc  <=~ dcache_s1_meta_clk_en & dcache_s2_req_no_alloc ;
             if ( dcache__GEN_63 )
                 begin 
                 end 
              else  
                 dcache_s2_uncached_resp_addr  <= dcache_uncachedResp_addr ; 
             dcache_s2_flush_valid_pre_tag_ecc  <= dcache_s1_flush_valid ;
             if ( dcache_s2_data_en ) 
                 dcache_s2_data  <=( dcache__s2_data_T_1 [0] ?  dcache_s2_data_s1_way_words_0_0 :32'h0)|( dcache__s2_data_T_1 [1] ?  dcache_s2_data_s1_way_words_1_0 :32'h0);
             if ( dcache_s1_valid_not_nacked ) 
                 dcache_s2_hit_way  <= dcache_s1_hit_way ;
             if ( dcache_s2_valid_cached_miss ) 
                 dcache_lrscAddr  <= dcache_s2_req_addr [31:6]; 
             dcache_s2_correct_REG  <= dcache_any_pstore_valid | dcache_s2_valid ;
             if ( dcache_s1_valid_not_nacked & dcache_s1_write )
                 begin  
                     dcache_pstore1_cmd  <= dcache_s1_req_cmd ; 
                     dcache_pstore1_addr  <= dcache_s1_vaddr ; 
                     dcache_pstore1_data  <= dcache_io_cpu_s1_data_data ; 
                     dcache_pstore1_way  <= dcache_s1_hit_way ; 
                     dcache_pstore1_mask  <= dcache_s1_mask ; 
                     dcache_pstore1_rmw_r  <= dcache__io_cpu_perf_canAcceptLoadThenLoad_T_1 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_2 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_3 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_29 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_31 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_32 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_33 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_34 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_38 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_39 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_40 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_41 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_42 |( dcache__io_cpu_perf_canAcceptLoadThenLoad_T_26 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_51 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_29 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_31 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_32 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_33 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_34 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_38 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_39 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_40 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_41 | dcache__io_cpu_perf_canAcceptLoadThenLoad_T_42 )& dcache__io_cpu_perf_canAcceptLoadThenLoad_T_51 ;
                 end  
             dcache_pstore_drain_on_miss_REG  <= dcache__io_cpu_s2_nack_output ;
             if ( dcache_advance_pstore1 )
                 begin  
                     dcache_pstore2_addr  <= dcache_pstore1_addr ; 
                     dcache_pstore2_way  <= dcache_pstore1_way ; 
                     dcache_pstore2_storegen_data_r  <= dcache_pstore1_storegen_data [7:0]; 
                     dcache_pstore2_storegen_data_r_1  <= dcache_pstore1_storegen_data [15:8]; 
                     dcache_pstore2_storegen_data_r_2  <= dcache_pstore1_storegen_data [23:16]; 
                     dcache_pstore2_storegen_data_r_3  <= dcache_pstore1_storegen_data [31:24]; 
                     dcache_pstore2_storegen_mask  <= dcache_pstore2_storegen_mask_mergedMask ;
                 end  
             dcache_io_cpu_s2_nack_cause_raw_REG  <= dcache_s1_raw_hazard ;
             if ( dcache__GEN_65 ) 
                 dcache_blockUncachedGrant  <=~ dcache_dataArb_grant_1 ;
              else  
                 dcache_blockUncachedGrant  <= dcache_dataArb_io_out_valid ; 
             dcache_s2_release_data_valid  <=1'h0; 
             dcache_io_cpu_s2_xcpt_REG  <= dcache_s1_xcpt_valid ;
             if ( dcache__io_cpu_replay_next_output ) 
                 dcache_s2_uncached_data_word  <= dcache_s1_uncached_data_word ; 
             dcache_doUncachedResp  <= dcache__io_cpu_replay_next_output ;
         end
    wire[1:0] dcache_tlb_pmp_io_prv;
    wire dcache_tlb_pmp_io_pmp_0_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_0_cfg_a;
    wire dcache_tlb_pmp_io_pmp_0_cfg_x;
    wire dcache_tlb_pmp_io_pmp_0_cfg_w;
    wire dcache_tlb_pmp_io_pmp_0_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_0_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_0_mask;
    wire dcache_tlb_pmp_io_pmp_1_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_1_cfg_a;
    wire dcache_tlb_pmp_io_pmp_1_cfg_x;
    wire dcache_tlb_pmp_io_pmp_1_cfg_w;
    wire dcache_tlb_pmp_io_pmp_1_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_1_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_1_mask;
    wire dcache_tlb_pmp_io_pmp_2_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_2_cfg_a;
    wire dcache_tlb_pmp_io_pmp_2_cfg_x;
    wire dcache_tlb_pmp_io_pmp_2_cfg_w;
    wire dcache_tlb_pmp_io_pmp_2_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_2_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_2_mask;
    wire dcache_tlb_pmp_io_pmp_3_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_3_cfg_a;
    wire dcache_tlb_pmp_io_pmp_3_cfg_x;
    wire dcache_tlb_pmp_io_pmp_3_cfg_w;
    wire dcache_tlb_pmp_io_pmp_3_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_3_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_3_mask;
    wire dcache_tlb_pmp_io_pmp_4_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_4_cfg_a;
    wire dcache_tlb_pmp_io_pmp_4_cfg_x;
    wire dcache_tlb_pmp_io_pmp_4_cfg_w;
    wire dcache_tlb_pmp_io_pmp_4_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_4_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_4_mask;
    wire dcache_tlb_pmp_io_pmp_5_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_5_cfg_a;
    wire dcache_tlb_pmp_io_pmp_5_cfg_x;
    wire dcache_tlb_pmp_io_pmp_5_cfg_w;
    wire dcache_tlb_pmp_io_pmp_5_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_5_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_5_mask;
    wire dcache_tlb_pmp_io_pmp_6_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_6_cfg_a;
    wire dcache_tlb_pmp_io_pmp_6_cfg_x;
    wire dcache_tlb_pmp_io_pmp_6_cfg_w;
    wire dcache_tlb_pmp_io_pmp_6_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_6_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_6_mask;
    wire dcache_tlb_pmp_io_pmp_7_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_7_cfg_a;
    wire dcache_tlb_pmp_io_pmp_7_cfg_x;
    wire dcache_tlb_pmp_io_pmp_7_cfg_w;
    wire dcache_tlb_pmp_io_pmp_7_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_7_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_7_mask;
    wire[31:0] dcache_tlb_pmp_io_addr;
    wire dcache_tlb_pmp_io_r;
    wire dcache_tlb_pmp_io_w;
    wire dcache_tlb_pmp_io_x;
    wire[1:0] dcache_pma_checker_pmp_io_prv;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_0_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_0_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_0_mask;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_1_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_1_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_1_mask;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_2_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_2_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_2_mask;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_3_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_3_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_3_mask;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_4_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_4_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_4_mask;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_5_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_5_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_5_mask;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_6_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_6_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_6_mask;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_7_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_7_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_7_mask;
    wire[31:0] dcache_pma_checker_pmp_io_addr;
    wire dcache_pma_checker_pmp_io_r;
    wire dcache_pma_checker_pmp_io_w;
    wire dcache_pma_checker_pmp_io_x;

    wire dcache_tlb_pmp_res_cur_cfg_l = dcache_tlb_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_cfg_a = dcache_tlb_pmp_io_pmp_7_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_addr = dcache_tlb_pmp_io_pmp_7_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_mask = dcache_tlb_pmp_io_pmp_7_mask ; 
    wire dcache_tlb_pmp_res_cur_1_cfg_l = dcache_tlb_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_1_cfg_a = dcache_tlb_pmp_io_pmp_6_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_1_addr = dcache_tlb_pmp_io_pmp_6_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_1_mask = dcache_tlb_pmp_io_pmp_6_mask ; 
    wire dcache_tlb_pmp_res_cur_2_cfg_l = dcache_tlb_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_2_cfg_a = dcache_tlb_pmp_io_pmp_5_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_2_addr = dcache_tlb_pmp_io_pmp_5_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_2_mask = dcache_tlb_pmp_io_pmp_5_mask ; 
    wire dcache_tlb_pmp_res_cur_3_cfg_l = dcache_tlb_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_3_cfg_a = dcache_tlb_pmp_io_pmp_4_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_3_addr = dcache_tlb_pmp_io_pmp_4_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_3_mask = dcache_tlb_pmp_io_pmp_4_mask ; 
    wire dcache_tlb_pmp_res_cur_4_cfg_l = dcache_tlb_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_4_cfg_a = dcache_tlb_pmp_io_pmp_3_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_4_addr = dcache_tlb_pmp_io_pmp_3_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_4_mask = dcache_tlb_pmp_io_pmp_3_mask ; 
    wire dcache_tlb_pmp_res_cur_5_cfg_l = dcache_tlb_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_5_cfg_a = dcache_tlb_pmp_io_pmp_2_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_5_addr = dcache_tlb_pmp_io_pmp_2_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_5_mask = dcache_tlb_pmp_io_pmp_2_mask ; 
    wire dcache_tlb_pmp_res_cur_6_cfg_l = dcache_tlb_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_6_cfg_a = dcache_tlb_pmp_io_pmp_1_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_6_addr = dcache_tlb_pmp_io_pmp_1_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_6_mask = dcache_tlb_pmp_io_pmp_1_mask ; 
    wire dcache_tlb_pmp_res_cur_7_cfg_l = dcache_tlb_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_7_cfg_a = dcache_tlb_pmp_io_pmp_0_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_7_addr = dcache_tlb_pmp_io_pmp_0_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_7_mask = dcache_tlb_pmp_io_pmp_0_mask ; 
    wire[1:0] dcache_tlb_pmp_pmp0_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_pmp0_cfg_a =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_1_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_2_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_3_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_4_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_5_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_6_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cur_7_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp_res_cfg_res =2'h0; 
    wire dcache_tlb_pmp_pmp0_cfg_l =1'h0; 
    wire[29:0] dcache_tlb_pmp_pmp0_addr =30'h0; 
    wire[31:0] dcache_tlb_pmp_pmp0_mask =32'h0; 
    wire dcache_tlb_pmp_default_0 = dcache_tlb_pmp_io_prv [1]; 
    wire dcache_tlb_pmp_pmp0_cfg_x = dcache_tlb_pmp_default_0 ; 
    wire dcache_tlb_pmp_pmp0_cfg_w = dcache_tlb_pmp_default_0 ; 
    wire dcache_tlb_pmp_pmp0_cfg_r = dcache_tlb_pmp_default_0 ; 
    wire dcache_tlb_pmp_res_hit = dcache_tlb_pmp_io_pmp_7_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_7_mask )==32'h0: dcache_tlb_pmp_io_pmp_7_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi ; 
  assign  dcache_tlb_pmp_res_hi = dcache_tlb_pmp__GEN ; 
    wire[1:0] dcache_tlb_pmp_res_hi_1 ; 
  assign  dcache_tlb_pmp_res_hi_1 = dcache_tlb_pmp__GEN ; 
    wire[1:0] dcache_tlb_pmp_res_hi_2 ; 
  assign  dcache_tlb_pmp_res_hi_2 = dcache_tlb_pmp__GEN ; 
    wire[1:0] dcache_tlb_pmp_res_hi_3 ; 
  assign  dcache_tlb_pmp_res_hi_3 = dcache_tlb_pmp__GEN ; 
    wire[1:0] dcache_tlb_pmp_res_hi_4 ; 
  assign  dcache_tlb_pmp_res_hi_4 = dcache_tlb_pmp__GEN ; 
    wire[1:0] dcache_tlb_pmp_res_hi_5 ; 
  assign  dcache_tlb_pmp_res_hi_5 = dcache_tlb_pmp__GEN ; 
    wire dcache_tlb_pmp_res_cur_cfg_r = dcache_tlb_pmp_io_pmp_7_cfg_r | dcache_tlb_pmp_res_ignore ; 
    wire dcache_tlb_pmp_res_cur_cfg_w = dcache_tlb_pmp_io_pmp_7_cfg_w | dcache_tlb_pmp_res_ignore ; 
    wire dcache_tlb_pmp_res_cur_cfg_x = dcache_tlb_pmp_io_pmp_7_cfg_x | dcache_tlb_pmp_res_ignore ; 
    wire dcache_tlb_pmp_res_hit_1 = dcache_tlb_pmp_io_pmp_6_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_6_mask )==32'h0: dcache_tlb_pmp_io_pmp_6_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_1 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_0 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_6 ; 
  assign  dcache_tlb_pmp_res_hi_6 = dcache_tlb_pmp__GEN_0 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_7 ; 
  assign  dcache_tlb_pmp_res_hi_7 = dcache_tlb_pmp__GEN_0 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_8 ; 
  assign  dcache_tlb_pmp_res_hi_8 = dcache_tlb_pmp__GEN_0 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_9 ; 
  assign  dcache_tlb_pmp_res_hi_9 = dcache_tlb_pmp__GEN_0 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_10 ; 
  assign  dcache_tlb_pmp_res_hi_10 = dcache_tlb_pmp__GEN_0 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_11 ; 
  assign  dcache_tlb_pmp_res_hi_11 = dcache_tlb_pmp__GEN_0 ; 
    wire dcache_tlb_pmp_res_cur_1_cfg_r = dcache_tlb_pmp_io_pmp_6_cfg_r | dcache_tlb_pmp_res_ignore_1 ; 
    wire dcache_tlb_pmp_res_cur_1_cfg_w = dcache_tlb_pmp_io_pmp_6_cfg_w | dcache_tlb_pmp_res_ignore_1 ; 
    wire dcache_tlb_pmp_res_cur_1_cfg_x = dcache_tlb_pmp_io_pmp_6_cfg_x | dcache_tlb_pmp_res_ignore_1 ; 
    wire dcache_tlb_pmp_res_hit_2 = dcache_tlb_pmp_io_pmp_5_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_5_mask )==32'h0: dcache_tlb_pmp_io_pmp_5_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_2 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_1 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_12 ; 
  assign  dcache_tlb_pmp_res_hi_12 = dcache_tlb_pmp__GEN_1 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_13 ; 
  assign  dcache_tlb_pmp_res_hi_13 = dcache_tlb_pmp__GEN_1 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_14 ; 
  assign  dcache_tlb_pmp_res_hi_14 = dcache_tlb_pmp__GEN_1 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_15 ; 
  assign  dcache_tlb_pmp_res_hi_15 = dcache_tlb_pmp__GEN_1 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_16 ; 
  assign  dcache_tlb_pmp_res_hi_16 = dcache_tlb_pmp__GEN_1 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_17 ; 
  assign  dcache_tlb_pmp_res_hi_17 = dcache_tlb_pmp__GEN_1 ; 
    wire dcache_tlb_pmp_res_cur_2_cfg_r = dcache_tlb_pmp_io_pmp_5_cfg_r | dcache_tlb_pmp_res_ignore_2 ; 
    wire dcache_tlb_pmp_res_cur_2_cfg_w = dcache_tlb_pmp_io_pmp_5_cfg_w | dcache_tlb_pmp_res_ignore_2 ; 
    wire dcache_tlb_pmp_res_cur_2_cfg_x = dcache_tlb_pmp_io_pmp_5_cfg_x | dcache_tlb_pmp_res_ignore_2 ; 
    wire dcache_tlb_pmp_res_hit_3 = dcache_tlb_pmp_io_pmp_4_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_4_mask )==32'h0: dcache_tlb_pmp_io_pmp_4_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_3 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_2 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_18 ; 
  assign  dcache_tlb_pmp_res_hi_18 = dcache_tlb_pmp__GEN_2 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_19 ; 
  assign  dcache_tlb_pmp_res_hi_19 = dcache_tlb_pmp__GEN_2 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_20 ; 
  assign  dcache_tlb_pmp_res_hi_20 = dcache_tlb_pmp__GEN_2 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_21 ; 
  assign  dcache_tlb_pmp_res_hi_21 = dcache_tlb_pmp__GEN_2 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_22 ; 
  assign  dcache_tlb_pmp_res_hi_22 = dcache_tlb_pmp__GEN_2 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_23 ; 
  assign  dcache_tlb_pmp_res_hi_23 = dcache_tlb_pmp__GEN_2 ; 
    wire dcache_tlb_pmp_res_cur_3_cfg_r = dcache_tlb_pmp_io_pmp_4_cfg_r | dcache_tlb_pmp_res_ignore_3 ; 
    wire dcache_tlb_pmp_res_cur_3_cfg_w = dcache_tlb_pmp_io_pmp_4_cfg_w | dcache_tlb_pmp_res_ignore_3 ; 
    wire dcache_tlb_pmp_res_cur_3_cfg_x = dcache_tlb_pmp_io_pmp_4_cfg_x | dcache_tlb_pmp_res_ignore_3 ; 
    wire dcache_tlb_pmp_res_hit_4 = dcache_tlb_pmp_io_pmp_3_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_3_mask )==32'h0: dcache_tlb_pmp_io_pmp_3_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_4 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_3 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_24 ; 
  assign  dcache_tlb_pmp_res_hi_24 = dcache_tlb_pmp__GEN_3 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_25 ; 
  assign  dcache_tlb_pmp_res_hi_25 = dcache_tlb_pmp__GEN_3 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_26 ; 
  assign  dcache_tlb_pmp_res_hi_26 = dcache_tlb_pmp__GEN_3 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_27 ; 
  assign  dcache_tlb_pmp_res_hi_27 = dcache_tlb_pmp__GEN_3 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_28 ; 
  assign  dcache_tlb_pmp_res_hi_28 = dcache_tlb_pmp__GEN_3 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_29 ; 
  assign  dcache_tlb_pmp_res_hi_29 = dcache_tlb_pmp__GEN_3 ; 
    wire dcache_tlb_pmp_res_cur_4_cfg_r = dcache_tlb_pmp_io_pmp_3_cfg_r | dcache_tlb_pmp_res_ignore_4 ; 
    wire dcache_tlb_pmp_res_cur_4_cfg_w = dcache_tlb_pmp_io_pmp_3_cfg_w | dcache_tlb_pmp_res_ignore_4 ; 
    wire dcache_tlb_pmp_res_cur_4_cfg_x = dcache_tlb_pmp_io_pmp_3_cfg_x | dcache_tlb_pmp_res_ignore_4 ; 
    wire dcache_tlb_pmp_res_hit_5 = dcache_tlb_pmp_io_pmp_2_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_2_mask )==32'h0: dcache_tlb_pmp_io_pmp_2_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_5 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_4 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_30 ; 
  assign  dcache_tlb_pmp_res_hi_30 = dcache_tlb_pmp__GEN_4 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_31 ; 
  assign  dcache_tlb_pmp_res_hi_31 = dcache_tlb_pmp__GEN_4 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_32 ; 
  assign  dcache_tlb_pmp_res_hi_32 = dcache_tlb_pmp__GEN_4 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_33 ; 
  assign  dcache_tlb_pmp_res_hi_33 = dcache_tlb_pmp__GEN_4 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_34 ; 
  assign  dcache_tlb_pmp_res_hi_34 = dcache_tlb_pmp__GEN_4 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_35 ; 
  assign  dcache_tlb_pmp_res_hi_35 = dcache_tlb_pmp__GEN_4 ; 
    wire dcache_tlb_pmp_res_cur_5_cfg_r = dcache_tlb_pmp_io_pmp_2_cfg_r | dcache_tlb_pmp_res_ignore_5 ; 
    wire dcache_tlb_pmp_res_cur_5_cfg_w = dcache_tlb_pmp_io_pmp_2_cfg_w | dcache_tlb_pmp_res_ignore_5 ; 
    wire dcache_tlb_pmp_res_cur_5_cfg_x = dcache_tlb_pmp_io_pmp_2_cfg_x | dcache_tlb_pmp_res_ignore_5 ; 
    wire dcache_tlb_pmp_res_hit_6 = dcache_tlb_pmp_io_pmp_1_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_1_mask )==32'h0: dcache_tlb_pmp_io_pmp_1_cfg_a [0]& dcache_tlb_pmp_io_addr >={ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_6 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_5 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_36 ; 
  assign  dcache_tlb_pmp_res_hi_36 = dcache_tlb_pmp__GEN_5 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_37 ; 
  assign  dcache_tlb_pmp_res_hi_37 = dcache_tlb_pmp__GEN_5 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_38 ; 
  assign  dcache_tlb_pmp_res_hi_38 = dcache_tlb_pmp__GEN_5 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_39 ; 
  assign  dcache_tlb_pmp_res_hi_39 = dcache_tlb_pmp__GEN_5 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_40 ; 
  assign  dcache_tlb_pmp_res_hi_40 = dcache_tlb_pmp__GEN_5 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_41 ; 
  assign  dcache_tlb_pmp_res_hi_41 = dcache_tlb_pmp__GEN_5 ; 
    wire dcache_tlb_pmp_res_cur_6_cfg_r = dcache_tlb_pmp_io_pmp_1_cfg_r | dcache_tlb_pmp_res_ignore_6 ; 
    wire dcache_tlb_pmp_res_cur_6_cfg_w = dcache_tlb_pmp_io_pmp_1_cfg_w | dcache_tlb_pmp_res_ignore_6 ; 
    wire dcache_tlb_pmp_res_cur_6_cfg_x = dcache_tlb_pmp_io_pmp_1_cfg_x | dcache_tlb_pmp_res_ignore_6 ; 
    wire dcache_tlb_pmp_res_hit_7 = dcache_tlb_pmp_io_pmp_0_cfg_a [1] ? (( dcache_tlb_pmp_io_addr ^{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0})&~ dcache_tlb_pmp_io_pmp_0_mask )==32'h0: dcache_tlb_pmp_io_pmp_0_cfg_a [0]& dcache_tlb_pmp_io_addr <{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}; 
    wire dcache_tlb_pmp_res_ignore_7 = dcache_tlb_pmp_default_0 &~ dcache_tlb_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] dcache_tlb_pmp__GEN_6 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_42 ; 
  assign  dcache_tlb_pmp_res_hi_42 = dcache_tlb_pmp__GEN_6 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_43 ; 
  assign  dcache_tlb_pmp_res_hi_43 = dcache_tlb_pmp__GEN_6 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_44 ; 
  assign  dcache_tlb_pmp_res_hi_44 = dcache_tlb_pmp__GEN_6 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_45 ; 
  assign  dcache_tlb_pmp_res_hi_45 = dcache_tlb_pmp__GEN_6 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_46 ; 
  assign  dcache_tlb_pmp_res_hi_46 = dcache_tlb_pmp__GEN_6 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_47 ; 
  assign  dcache_tlb_pmp_res_hi_47 = dcache_tlb_pmp__GEN_6 ; 
    wire dcache_tlb_pmp_res_cur_7_cfg_r = dcache_tlb_pmp_io_pmp_0_cfg_r | dcache_tlb_pmp_res_ignore_7 ; 
    wire dcache_tlb_pmp_res_cur_7_cfg_w = dcache_tlb_pmp_io_pmp_0_cfg_w | dcache_tlb_pmp_res_ignore_7 ; 
    wire dcache_tlb_pmp_res_cur_7_cfg_x = dcache_tlb_pmp_io_pmp_0_cfg_x | dcache_tlb_pmp_res_ignore_7 ; 
    wire dcache_tlb_pmp_res_cfg_l = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_l : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_l : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_l : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_l : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_l : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_l : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_l : dcache_tlb_pmp_res_hit & dcache_tlb_pmp_res_cur_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cfg_a = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_a : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_a : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_a : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_a : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_a : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_a : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_a : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_a :2'h0; 
    wire dcache_tlb_pmp_res_cfg_x = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_x : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_x : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_x : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_x : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_x : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_x : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_x : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_x : dcache_tlb_pmp_pmp0_cfg_x ; 
    wire dcache_tlb_pmp_res_cfg_w = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_w : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_w : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_w : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_w : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_w : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_w : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_w : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_w : dcache_tlb_pmp_pmp0_cfg_w ; 
    wire dcache_tlb_pmp_res_cfg_r = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_r : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_r : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_r : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_r : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_r : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_r : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_r : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_r : dcache_tlb_pmp_pmp0_cfg_r ; 
    wire[29:0] dcache_tlb_pmp_res_addr = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_addr : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_addr : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_addr : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_addr : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_addr : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_addr : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_addr : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_addr :30'h0; 
    wire[31:0] dcache_tlb_pmp_res_mask = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_mask : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_mask : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_mask : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_mask : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_mask : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_mask : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_mask : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_mask :32'h0; 
  assign  dcache_tlb_pmp_io_r = dcache_tlb_pmp_res_cfg_r ; 
  assign  dcache_tlb_pmp_io_w = dcache_tlb_pmp_res_cfg_w ; 
  assign  dcache_tlb_pmp_io_x = dcache_tlb_pmp_res_cfg_x ;
      
    wire dcache_tlb_entries_barrier_io_x_u;
    wire dcache_tlb_entries_barrier_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_io_x_ae_final;
    wire dcache_tlb_entries_barrier_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_io_x_pf;
    wire dcache_tlb_entries_barrier_io_x_gf;
    wire dcache_tlb_entries_barrier_io_x_sw;
    wire dcache_tlb_entries_barrier_io_x_sx;
    wire dcache_tlb_entries_barrier_io_x_sr;
    wire dcache_tlb_entries_barrier_io_x_hw;
    wire dcache_tlb_entries_barrier_io_x_hx;
    wire dcache_tlb_entries_barrier_io_x_hr;
    wire dcache_tlb_entries_barrier_io_x_pw;
    wire dcache_tlb_entries_barrier_io_x_px;
    wire dcache_tlb_entries_barrier_io_x_pr;
    wire dcache_tlb_entries_barrier_io_x_ppp;
    wire dcache_tlb_entries_barrier_io_x_pal;
    wire dcache_tlb_entries_barrier_io_x_paa;
    wire dcache_tlb_entries_barrier_io_x_eff;
    wire dcache_tlb_entries_barrier_io_x_c;
    wire dcache_tlb_entries_barrier_io_y_u;
    wire dcache_tlb_entries_barrier_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_io_y_ae_final;
    wire dcache_tlb_entries_barrier_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_io_y_pf;
    wire dcache_tlb_entries_barrier_io_y_gf;
    wire dcache_tlb_entries_barrier_io_y_sw;
    wire dcache_tlb_entries_barrier_io_y_sx;
    wire dcache_tlb_entries_barrier_io_y_sr;
    wire dcache_tlb_entries_barrier_io_y_hw;
    wire dcache_tlb_entries_barrier_io_y_hx;
    wire dcache_tlb_entries_barrier_io_y_hr;
    wire dcache_tlb_entries_barrier_io_y_pw;
    wire dcache_tlb_entries_barrier_io_y_px;
    wire dcache_tlb_entries_barrier_io_y_pr;
    wire dcache_tlb_entries_barrier_io_y_ppp;
    wire dcache_tlb_entries_barrier_io_y_pal;
    wire dcache_tlb_entries_barrier_io_y_paa;
    wire dcache_tlb_entries_barrier_io_y_eff;
    wire dcache_tlb_entries_barrier_io_y_c;
    wire dcache_tlb_entries_barrier_1_io_x_u;
    wire dcache_tlb_entries_barrier_1_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_1_io_x_ae_final;
    wire dcache_tlb_entries_barrier_1_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_1_io_x_pf;
    wire dcache_tlb_entries_barrier_1_io_x_gf;
    wire dcache_tlb_entries_barrier_1_io_x_sw;
    wire dcache_tlb_entries_barrier_1_io_x_sx;
    wire dcache_tlb_entries_barrier_1_io_x_sr;
    wire dcache_tlb_entries_barrier_1_io_x_hw;
    wire dcache_tlb_entries_barrier_1_io_x_hx;
    wire dcache_tlb_entries_barrier_1_io_x_hr;
    wire dcache_tlb_entries_barrier_1_io_x_pw;
    wire dcache_tlb_entries_barrier_1_io_x_px;
    wire dcache_tlb_entries_barrier_1_io_x_pr;
    wire dcache_tlb_entries_barrier_1_io_x_ppp;
    wire dcache_tlb_entries_barrier_1_io_x_pal;
    wire dcache_tlb_entries_barrier_1_io_x_paa;
    wire dcache_tlb_entries_barrier_1_io_x_eff;
    wire dcache_tlb_entries_barrier_1_io_x_c;
    wire dcache_tlb_entries_barrier_1_io_y_u;
    wire dcache_tlb_entries_barrier_1_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_1_io_y_ae_final;
    wire dcache_tlb_entries_barrier_1_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_1_io_y_pf;
    wire dcache_tlb_entries_barrier_1_io_y_gf;
    wire dcache_tlb_entries_barrier_1_io_y_sw;
    wire dcache_tlb_entries_barrier_1_io_y_sx;
    wire dcache_tlb_entries_barrier_1_io_y_sr;
    wire dcache_tlb_entries_barrier_1_io_y_hw;
    wire dcache_tlb_entries_barrier_1_io_y_hx;
    wire dcache_tlb_entries_barrier_1_io_y_hr;
    wire dcache_tlb_entries_barrier_1_io_y_pw;
    wire dcache_tlb_entries_barrier_1_io_y_px;
    wire dcache_tlb_entries_barrier_1_io_y_pr;
    wire dcache_tlb_entries_barrier_1_io_y_ppp;
    wire dcache_tlb_entries_barrier_1_io_y_pal;
    wire dcache_tlb_entries_barrier_1_io_y_paa;
    wire dcache_tlb_entries_barrier_1_io_y_eff;
    wire dcache_tlb_entries_barrier_1_io_y_c;
    wire dcache_tlb_entries_barrier_2_io_x_u;
    wire dcache_tlb_entries_barrier_2_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_2_io_x_ae_final;
    wire dcache_tlb_entries_barrier_2_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_2_io_x_pf;
    wire dcache_tlb_entries_barrier_2_io_x_gf;
    wire dcache_tlb_entries_barrier_2_io_x_sw;
    wire dcache_tlb_entries_barrier_2_io_x_sx;
    wire dcache_tlb_entries_barrier_2_io_x_sr;
    wire dcache_tlb_entries_barrier_2_io_x_hw;
    wire dcache_tlb_entries_barrier_2_io_x_hx;
    wire dcache_tlb_entries_barrier_2_io_x_hr;
    wire dcache_tlb_entries_barrier_2_io_x_pw;
    wire dcache_tlb_entries_barrier_2_io_x_px;
    wire dcache_tlb_entries_barrier_2_io_x_pr;
    wire dcache_tlb_entries_barrier_2_io_x_ppp;
    wire dcache_tlb_entries_barrier_2_io_x_pal;
    wire dcache_tlb_entries_barrier_2_io_x_paa;
    wire dcache_tlb_entries_barrier_2_io_x_eff;
    wire dcache_tlb_entries_barrier_2_io_x_c;
    wire dcache_tlb_entries_barrier_2_io_y_u;
    wire dcache_tlb_entries_barrier_2_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_2_io_y_ae_final;
    wire dcache_tlb_entries_barrier_2_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_2_io_y_pf;
    wire dcache_tlb_entries_barrier_2_io_y_gf;
    wire dcache_tlb_entries_barrier_2_io_y_sw;
    wire dcache_tlb_entries_barrier_2_io_y_sx;
    wire dcache_tlb_entries_barrier_2_io_y_sr;
    wire dcache_tlb_entries_barrier_2_io_y_hw;
    wire dcache_tlb_entries_barrier_2_io_y_hx;
    wire dcache_tlb_entries_barrier_2_io_y_hr;
    wire dcache_tlb_entries_barrier_2_io_y_pw;
    wire dcache_tlb_entries_barrier_2_io_y_px;
    wire dcache_tlb_entries_barrier_2_io_y_pr;
    wire dcache_tlb_entries_barrier_2_io_y_ppp;
    wire dcache_tlb_entries_barrier_2_io_y_pal;
    wire dcache_tlb_entries_barrier_2_io_y_paa;
    wire dcache_tlb_entries_barrier_2_io_y_eff;
    wire dcache_tlb_entries_barrier_2_io_y_c;
    wire dcache_tlb_entries_barrier_3_io_x_u;
    wire dcache_tlb_entries_barrier_3_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_3_io_x_ae_final;
    wire dcache_tlb_entries_barrier_3_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_3_io_x_pf;
    wire dcache_tlb_entries_barrier_3_io_x_gf;
    wire dcache_tlb_entries_barrier_3_io_x_sw;
    wire dcache_tlb_entries_barrier_3_io_x_sx;
    wire dcache_tlb_entries_barrier_3_io_x_sr;
    wire dcache_tlb_entries_barrier_3_io_x_hw;
    wire dcache_tlb_entries_barrier_3_io_x_hx;
    wire dcache_tlb_entries_barrier_3_io_x_hr;
    wire dcache_tlb_entries_barrier_3_io_x_pw;
    wire dcache_tlb_entries_barrier_3_io_x_px;
    wire dcache_tlb_entries_barrier_3_io_x_pr;
    wire dcache_tlb_entries_barrier_3_io_x_ppp;
    wire dcache_tlb_entries_barrier_3_io_x_pal;
    wire dcache_tlb_entries_barrier_3_io_x_paa;
    wire dcache_tlb_entries_barrier_3_io_x_eff;
    wire dcache_tlb_entries_barrier_3_io_x_c;
    wire dcache_tlb_entries_barrier_3_io_y_u;
    wire dcache_tlb_entries_barrier_3_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_3_io_y_ae_final;
    wire dcache_tlb_entries_barrier_3_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_3_io_y_pf;
    wire dcache_tlb_entries_barrier_3_io_y_gf;
    wire dcache_tlb_entries_barrier_3_io_y_sw;
    wire dcache_tlb_entries_barrier_3_io_y_sx;
    wire dcache_tlb_entries_barrier_3_io_y_sr;
    wire dcache_tlb_entries_barrier_3_io_y_hw;
    wire dcache_tlb_entries_barrier_3_io_y_hx;
    wire dcache_tlb_entries_barrier_3_io_y_hr;
    wire dcache_tlb_entries_barrier_3_io_y_pw;
    wire dcache_tlb_entries_barrier_3_io_y_px;
    wire dcache_tlb_entries_barrier_3_io_y_pr;
    wire dcache_tlb_entries_barrier_3_io_y_ppp;
    wire dcache_tlb_entries_barrier_3_io_y_pal;
    wire dcache_tlb_entries_barrier_3_io_y_paa;
    wire dcache_tlb_entries_barrier_3_io_y_eff;
    wire dcache_tlb_entries_barrier_3_io_y_c;
    wire dcache_tlb_entries_barrier_4_io_x_u;
    wire dcache_tlb_entries_barrier_4_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_4_io_x_ae_final;
    wire dcache_tlb_entries_barrier_4_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_4_io_x_pf;
    wire dcache_tlb_entries_barrier_4_io_x_gf;
    wire dcache_tlb_entries_barrier_4_io_x_sw;
    wire dcache_tlb_entries_barrier_4_io_x_sx;
    wire dcache_tlb_entries_barrier_4_io_x_sr;
    wire dcache_tlb_entries_barrier_4_io_x_hw;
    wire dcache_tlb_entries_barrier_4_io_x_hx;
    wire dcache_tlb_entries_barrier_4_io_x_hr;
    wire dcache_tlb_entries_barrier_4_io_x_pw;
    wire dcache_tlb_entries_barrier_4_io_x_px;
    wire dcache_tlb_entries_barrier_4_io_x_pr;
    wire dcache_tlb_entries_barrier_4_io_x_ppp;
    wire dcache_tlb_entries_barrier_4_io_x_pal;
    wire dcache_tlb_entries_barrier_4_io_x_paa;
    wire dcache_tlb_entries_barrier_4_io_x_eff;
    wire dcache_tlb_entries_barrier_4_io_x_c;
    wire dcache_tlb_entries_barrier_4_io_y_u;
    wire dcache_tlb_entries_barrier_4_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_4_io_y_ae_final;
    wire dcache_tlb_entries_barrier_4_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_4_io_y_pf;
    wire dcache_tlb_entries_barrier_4_io_y_gf;
    wire dcache_tlb_entries_barrier_4_io_y_sw;
    wire dcache_tlb_entries_barrier_4_io_y_sx;
    wire dcache_tlb_entries_barrier_4_io_y_sr;
    wire dcache_tlb_entries_barrier_4_io_y_hw;
    wire dcache_tlb_entries_barrier_4_io_y_hx;
    wire dcache_tlb_entries_barrier_4_io_y_hr;
    wire dcache_tlb_entries_barrier_4_io_y_pw;
    wire dcache_tlb_entries_barrier_4_io_y_px;
    wire dcache_tlb_entries_barrier_4_io_y_pr;
    wire dcache_tlb_entries_barrier_4_io_y_ppp;
    wire dcache_tlb_entries_barrier_4_io_y_pal;
    wire dcache_tlb_entries_barrier_4_io_y_paa;
    wire dcache_tlb_entries_barrier_4_io_y_eff;
    wire dcache_tlb_entries_barrier_4_io_y_c;
    wire dcache_tlb_entries_barrier_5_io_x_u;
    wire dcache_tlb_entries_barrier_5_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_5_io_x_ae_final;
    wire dcache_tlb_entries_barrier_5_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_5_io_x_pf;
    wire dcache_tlb_entries_barrier_5_io_x_gf;
    wire dcache_tlb_entries_barrier_5_io_x_sw;
    wire dcache_tlb_entries_barrier_5_io_x_sx;
    wire dcache_tlb_entries_barrier_5_io_x_sr;
    wire dcache_tlb_entries_barrier_5_io_x_hw;
    wire dcache_tlb_entries_barrier_5_io_x_hx;
    wire dcache_tlb_entries_barrier_5_io_x_hr;
    wire dcache_tlb_entries_barrier_5_io_x_pw;
    wire dcache_tlb_entries_barrier_5_io_x_px;
    wire dcache_tlb_entries_barrier_5_io_x_pr;
    wire dcache_tlb_entries_barrier_5_io_x_ppp;
    wire dcache_tlb_entries_barrier_5_io_x_pal;
    wire dcache_tlb_entries_barrier_5_io_x_paa;
    wire dcache_tlb_entries_barrier_5_io_x_eff;
    wire dcache_tlb_entries_barrier_5_io_x_c;
    wire dcache_tlb_entries_barrier_5_io_y_u;
    wire dcache_tlb_entries_barrier_5_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_5_io_y_ae_final;
    wire dcache_tlb_entries_barrier_5_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_5_io_y_pf;
    wire dcache_tlb_entries_barrier_5_io_y_gf;
    wire dcache_tlb_entries_barrier_5_io_y_sw;
    wire dcache_tlb_entries_barrier_5_io_y_sx;
    wire dcache_tlb_entries_barrier_5_io_y_sr;
    wire dcache_tlb_entries_barrier_5_io_y_hw;
    wire dcache_tlb_entries_barrier_5_io_y_hx;
    wire dcache_tlb_entries_barrier_5_io_y_hr;
    wire dcache_tlb_entries_barrier_5_io_y_pw;
    wire dcache_tlb_entries_barrier_5_io_y_px;
    wire dcache_tlb_entries_barrier_5_io_y_pr;
    wire dcache_tlb_entries_barrier_5_io_y_ppp;
    wire dcache_tlb_entries_barrier_5_io_y_pal;
    wire dcache_tlb_entries_barrier_5_io_y_paa;
    wire dcache_tlb_entries_barrier_5_io_y_eff;
    wire dcache_tlb_entries_barrier_5_io_y_c;
    wire dcache_pma_checker_entries_barrier_io_x_u;
    wire dcache_pma_checker_entries_barrier_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_io_x_pf;
    wire dcache_pma_checker_entries_barrier_io_x_gf;
    wire dcache_pma_checker_entries_barrier_io_x_sw;
    wire dcache_pma_checker_entries_barrier_io_x_sx;
    wire dcache_pma_checker_entries_barrier_io_x_sr;
    wire dcache_pma_checker_entries_barrier_io_x_hw;
    wire dcache_pma_checker_entries_barrier_io_x_hx;
    wire dcache_pma_checker_entries_barrier_io_x_hr;
    wire dcache_pma_checker_entries_barrier_io_x_pw;
    wire dcache_pma_checker_entries_barrier_io_x_px;
    wire dcache_pma_checker_entries_barrier_io_x_pr;
    wire dcache_pma_checker_entries_barrier_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_io_x_pal;
    wire dcache_pma_checker_entries_barrier_io_x_paa;
    wire dcache_pma_checker_entries_barrier_io_x_eff;
    wire dcache_pma_checker_entries_barrier_io_x_c;
    wire dcache_pma_checker_entries_barrier_io_y_u;
    wire dcache_pma_checker_entries_barrier_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_io_y_pf;
    wire dcache_pma_checker_entries_barrier_io_y_gf;
    wire dcache_pma_checker_entries_barrier_io_y_sw;
    wire dcache_pma_checker_entries_barrier_io_y_sx;
    wire dcache_pma_checker_entries_barrier_io_y_sr;
    wire dcache_pma_checker_entries_barrier_io_y_hw;
    wire dcache_pma_checker_entries_barrier_io_y_hx;
    wire dcache_pma_checker_entries_barrier_io_y_hr;
    wire dcache_pma_checker_entries_barrier_io_y_pw;
    wire dcache_pma_checker_entries_barrier_io_y_px;
    wire dcache_pma_checker_entries_barrier_io_y_pr;
    wire dcache_pma_checker_entries_barrier_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_io_y_pal;
    wire dcache_pma_checker_entries_barrier_io_y_paa;
    wire dcache_pma_checker_entries_barrier_io_y_eff;
    wire dcache_pma_checker_entries_barrier_io_y_c;
    wire dcache_pma_checker_entries_barrier_1_io_x_u;
    wire dcache_pma_checker_entries_barrier_1_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_1_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_1_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_1_io_x_pf;
    wire dcache_pma_checker_entries_barrier_1_io_x_gf;
    wire dcache_pma_checker_entries_barrier_1_io_x_sw;
    wire dcache_pma_checker_entries_barrier_1_io_x_sx;
    wire dcache_pma_checker_entries_barrier_1_io_x_sr;
    wire dcache_pma_checker_entries_barrier_1_io_x_hw;
    wire dcache_pma_checker_entries_barrier_1_io_x_hx;
    wire dcache_pma_checker_entries_barrier_1_io_x_hr;
    wire dcache_pma_checker_entries_barrier_1_io_x_pw;
    wire dcache_pma_checker_entries_barrier_1_io_x_px;
    wire dcache_pma_checker_entries_barrier_1_io_x_pr;
    wire dcache_pma_checker_entries_barrier_1_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_1_io_x_pal;
    wire dcache_pma_checker_entries_barrier_1_io_x_paa;
    wire dcache_pma_checker_entries_barrier_1_io_x_eff;
    wire dcache_pma_checker_entries_barrier_1_io_x_c;
    wire dcache_pma_checker_entries_barrier_1_io_y_u;
    wire dcache_pma_checker_entries_barrier_1_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_1_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_1_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_1_io_y_pf;
    wire dcache_pma_checker_entries_barrier_1_io_y_gf;
    wire dcache_pma_checker_entries_barrier_1_io_y_sw;
    wire dcache_pma_checker_entries_barrier_1_io_y_sx;
    wire dcache_pma_checker_entries_barrier_1_io_y_sr;
    wire dcache_pma_checker_entries_barrier_1_io_y_hw;
    wire dcache_pma_checker_entries_barrier_1_io_y_hx;
    wire dcache_pma_checker_entries_barrier_1_io_y_hr;
    wire dcache_pma_checker_entries_barrier_1_io_y_pw;
    wire dcache_pma_checker_entries_barrier_1_io_y_px;
    wire dcache_pma_checker_entries_barrier_1_io_y_pr;
    wire dcache_pma_checker_entries_barrier_1_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_1_io_y_pal;
    wire dcache_pma_checker_entries_barrier_1_io_y_paa;
    wire dcache_pma_checker_entries_barrier_1_io_y_eff;
    wire dcache_pma_checker_entries_barrier_1_io_y_c;
    wire dcache_pma_checker_entries_barrier_2_io_x_u;
    wire dcache_pma_checker_entries_barrier_2_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_2_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_2_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_2_io_x_pf;
    wire dcache_pma_checker_entries_barrier_2_io_x_gf;
    wire dcache_pma_checker_entries_barrier_2_io_x_sw;
    wire dcache_pma_checker_entries_barrier_2_io_x_sx;
    wire dcache_pma_checker_entries_barrier_2_io_x_sr;
    wire dcache_pma_checker_entries_barrier_2_io_x_hw;
    wire dcache_pma_checker_entries_barrier_2_io_x_hx;
    wire dcache_pma_checker_entries_barrier_2_io_x_hr;
    wire dcache_pma_checker_entries_barrier_2_io_x_pw;
    wire dcache_pma_checker_entries_barrier_2_io_x_px;
    wire dcache_pma_checker_entries_barrier_2_io_x_pr;
    wire dcache_pma_checker_entries_barrier_2_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_2_io_x_pal;
    wire dcache_pma_checker_entries_barrier_2_io_x_paa;
    wire dcache_pma_checker_entries_barrier_2_io_x_eff;
    wire dcache_pma_checker_entries_barrier_2_io_x_c;
    wire dcache_pma_checker_entries_barrier_2_io_y_u;
    wire dcache_pma_checker_entries_barrier_2_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_2_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_2_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_2_io_y_pf;
    wire dcache_pma_checker_entries_barrier_2_io_y_gf;
    wire dcache_pma_checker_entries_barrier_2_io_y_sw;
    wire dcache_pma_checker_entries_barrier_2_io_y_sx;
    wire dcache_pma_checker_entries_barrier_2_io_y_sr;
    wire dcache_pma_checker_entries_barrier_2_io_y_hw;
    wire dcache_pma_checker_entries_barrier_2_io_y_hx;
    wire dcache_pma_checker_entries_barrier_2_io_y_hr;
    wire dcache_pma_checker_entries_barrier_2_io_y_pw;
    wire dcache_pma_checker_entries_barrier_2_io_y_px;
    wire dcache_pma_checker_entries_barrier_2_io_y_pr;
    wire dcache_pma_checker_entries_barrier_2_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_2_io_y_pal;
    wire dcache_pma_checker_entries_barrier_2_io_y_paa;
    wire dcache_pma_checker_entries_barrier_2_io_y_eff;
    wire dcache_pma_checker_entries_barrier_2_io_y_c;
    wire dcache_pma_checker_entries_barrier_3_io_x_u;
    wire dcache_pma_checker_entries_barrier_3_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_3_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_3_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_3_io_x_pf;
    wire dcache_pma_checker_entries_barrier_3_io_x_gf;
    wire dcache_pma_checker_entries_barrier_3_io_x_sw;
    wire dcache_pma_checker_entries_barrier_3_io_x_sx;
    wire dcache_pma_checker_entries_barrier_3_io_x_sr;
    wire dcache_pma_checker_entries_barrier_3_io_x_hw;
    wire dcache_pma_checker_entries_barrier_3_io_x_hx;
    wire dcache_pma_checker_entries_barrier_3_io_x_hr;
    wire dcache_pma_checker_entries_barrier_3_io_x_pw;
    wire dcache_pma_checker_entries_barrier_3_io_x_px;
    wire dcache_pma_checker_entries_barrier_3_io_x_pr;
    wire dcache_pma_checker_entries_barrier_3_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_3_io_x_pal;
    wire dcache_pma_checker_entries_barrier_3_io_x_paa;
    wire dcache_pma_checker_entries_barrier_3_io_x_eff;
    wire dcache_pma_checker_entries_barrier_3_io_x_c;
    wire dcache_pma_checker_entries_barrier_3_io_y_u;
    wire dcache_pma_checker_entries_barrier_3_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_3_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_3_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_3_io_y_pf;
    wire dcache_pma_checker_entries_barrier_3_io_y_gf;
    wire dcache_pma_checker_entries_barrier_3_io_y_sw;
    wire dcache_pma_checker_entries_barrier_3_io_y_sx;
    wire dcache_pma_checker_entries_barrier_3_io_y_sr;
    wire dcache_pma_checker_entries_barrier_3_io_y_hw;
    wire dcache_pma_checker_entries_barrier_3_io_y_hx;
    wire dcache_pma_checker_entries_barrier_3_io_y_hr;
    wire dcache_pma_checker_entries_barrier_3_io_y_pw;
    wire dcache_pma_checker_entries_barrier_3_io_y_px;
    wire dcache_pma_checker_entries_barrier_3_io_y_pr;
    wire dcache_pma_checker_entries_barrier_3_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_3_io_y_pal;
    wire dcache_pma_checker_entries_barrier_3_io_y_paa;
    wire dcache_pma_checker_entries_barrier_3_io_y_eff;
    wire dcache_pma_checker_entries_barrier_3_io_y_c;
    wire dcache_pma_checker_entries_barrier_4_io_x_u;
    wire dcache_pma_checker_entries_barrier_4_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_4_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_4_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_4_io_x_pf;
    wire dcache_pma_checker_entries_barrier_4_io_x_gf;
    wire dcache_pma_checker_entries_barrier_4_io_x_sw;
    wire dcache_pma_checker_entries_barrier_4_io_x_sx;
    wire dcache_pma_checker_entries_barrier_4_io_x_sr;
    wire dcache_pma_checker_entries_barrier_4_io_x_hw;
    wire dcache_pma_checker_entries_barrier_4_io_x_hx;
    wire dcache_pma_checker_entries_barrier_4_io_x_hr;
    wire dcache_pma_checker_entries_barrier_4_io_x_pw;
    wire dcache_pma_checker_entries_barrier_4_io_x_px;
    wire dcache_pma_checker_entries_barrier_4_io_x_pr;
    wire dcache_pma_checker_entries_barrier_4_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_4_io_x_pal;
    wire dcache_pma_checker_entries_barrier_4_io_x_paa;
    wire dcache_pma_checker_entries_barrier_4_io_x_eff;
    wire dcache_pma_checker_entries_barrier_4_io_x_c;
    wire dcache_pma_checker_entries_barrier_4_io_y_u;
    wire dcache_pma_checker_entries_barrier_4_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_4_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_4_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_4_io_y_pf;
    wire dcache_pma_checker_entries_barrier_4_io_y_gf;
    wire dcache_pma_checker_entries_barrier_4_io_y_sw;
    wire dcache_pma_checker_entries_barrier_4_io_y_sx;
    wire dcache_pma_checker_entries_barrier_4_io_y_sr;
    wire dcache_pma_checker_entries_barrier_4_io_y_hw;
    wire dcache_pma_checker_entries_barrier_4_io_y_hx;
    wire dcache_pma_checker_entries_barrier_4_io_y_hr;
    wire dcache_pma_checker_entries_barrier_4_io_y_pw;
    wire dcache_pma_checker_entries_barrier_4_io_y_px;
    wire dcache_pma_checker_entries_barrier_4_io_y_pr;
    wire dcache_pma_checker_entries_barrier_4_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_4_io_y_pal;
    wire dcache_pma_checker_entries_barrier_4_io_y_paa;
    wire dcache_pma_checker_entries_barrier_4_io_y_eff;
    wire dcache_pma_checker_entries_barrier_4_io_y_c;
    wire dcache_pma_checker_entries_barrier_5_io_x_u;
    wire dcache_pma_checker_entries_barrier_5_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_5_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_5_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_5_io_x_pf;
    wire dcache_pma_checker_entries_barrier_5_io_x_gf;
    wire dcache_pma_checker_entries_barrier_5_io_x_sw;
    wire dcache_pma_checker_entries_barrier_5_io_x_sx;
    wire dcache_pma_checker_entries_barrier_5_io_x_sr;
    wire dcache_pma_checker_entries_barrier_5_io_x_hw;
    wire dcache_pma_checker_entries_barrier_5_io_x_hx;
    wire dcache_pma_checker_entries_barrier_5_io_x_hr;
    wire dcache_pma_checker_entries_barrier_5_io_x_pw;
    wire dcache_pma_checker_entries_barrier_5_io_x_px;
    wire dcache_pma_checker_entries_barrier_5_io_x_pr;
    wire dcache_pma_checker_entries_barrier_5_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_5_io_x_pal;
    wire dcache_pma_checker_entries_barrier_5_io_x_paa;
    wire dcache_pma_checker_entries_barrier_5_io_x_eff;
    wire dcache_pma_checker_entries_barrier_5_io_x_c;
    wire dcache_pma_checker_entries_barrier_5_io_y_u;
    wire dcache_pma_checker_entries_barrier_5_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_5_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_5_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_5_io_y_pf;
    wire dcache_pma_checker_entries_barrier_5_io_y_gf;
    wire dcache_pma_checker_entries_barrier_5_io_y_sw;
    wire dcache_pma_checker_entries_barrier_5_io_y_sx;
    wire dcache_pma_checker_entries_barrier_5_io_y_sr;
    wire dcache_pma_checker_entries_barrier_5_io_y_hw;
    wire dcache_pma_checker_entries_barrier_5_io_y_hx;
    wire dcache_pma_checker_entries_barrier_5_io_y_hr;
    wire dcache_pma_checker_entries_barrier_5_io_y_pw;
    wire dcache_pma_checker_entries_barrier_5_io_y_px;
    wire dcache_pma_checker_entries_barrier_5_io_y_pr;
    wire dcache_pma_checker_entries_barrier_5_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_5_io_y_pal;
    wire dcache_pma_checker_entries_barrier_5_io_y_paa;
    wire dcache_pma_checker_entries_barrier_5_io_y_eff;
    wire dcache_pma_checker_entries_barrier_5_io_y_c;

    assign  dcache_tlb_entries_barrier_io_y_u = dcache_tlb_entries_barrier_io_x_u ; 
  assign  dcache_tlb_entries_barrier_io_y_ae_ptw = dcache_tlb_entries_barrier_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_io_y_ae_final = dcache_tlb_entries_barrier_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_io_y_ae_stage2 = dcache_tlb_entries_barrier_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_io_y_pf = dcache_tlb_entries_barrier_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_io_y_gf = dcache_tlb_entries_barrier_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_io_y_sw = dcache_tlb_entries_barrier_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_io_y_sx = dcache_tlb_entries_barrier_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_io_y_sr = dcache_tlb_entries_barrier_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_io_y_hw = dcache_tlb_entries_barrier_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_io_y_hx = dcache_tlb_entries_barrier_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_io_y_hr = dcache_tlb_entries_barrier_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_io_y_pw = dcache_tlb_entries_barrier_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_io_y_px = dcache_tlb_entries_barrier_io_x_px ; 
  assign  dcache_tlb_entries_barrier_io_y_pr = dcache_tlb_entries_barrier_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_io_y_ppp = dcache_tlb_entries_barrier_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_io_y_pal = dcache_tlb_entries_barrier_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_io_y_paa = dcache_tlb_entries_barrier_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_io_y_eff = dcache_tlb_entries_barrier_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_io_y_c = dcache_tlb_entries_barrier_io_x_c ;
    assign  dcache_tlb_entries_barrier_1_io_y_u = dcache_tlb_entries_barrier_1_io_x_u ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ae_ptw = dcache_tlb_entries_barrier_1_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ae_final = dcache_tlb_entries_barrier_1_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ae_stage2 = dcache_tlb_entries_barrier_1_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pf = dcache_tlb_entries_barrier_1_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_1_io_y_gf = dcache_tlb_entries_barrier_1_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_1_io_y_sw = dcache_tlb_entries_barrier_1_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_sx = dcache_tlb_entries_barrier_1_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_1_io_y_sr = dcache_tlb_entries_barrier_1_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_1_io_y_hw = dcache_tlb_entries_barrier_1_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_hx = dcache_tlb_entries_barrier_1_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_1_io_y_hr = dcache_tlb_entries_barrier_1_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pw = dcache_tlb_entries_barrier_1_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_px = dcache_tlb_entries_barrier_1_io_x_px ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pr = dcache_tlb_entries_barrier_1_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ppp = dcache_tlb_entries_barrier_1_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pal = dcache_tlb_entries_barrier_1_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_1_io_y_paa = dcache_tlb_entries_barrier_1_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_1_io_y_eff = dcache_tlb_entries_barrier_1_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_1_io_y_c = dcache_tlb_entries_barrier_1_io_x_c ;
    assign  dcache_tlb_entries_barrier_2_io_y_u = dcache_tlb_entries_barrier_2_io_x_u ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ae_ptw = dcache_tlb_entries_barrier_2_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ae_final = dcache_tlb_entries_barrier_2_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ae_stage2 = dcache_tlb_entries_barrier_2_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pf = dcache_tlb_entries_barrier_2_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_2_io_y_gf = dcache_tlb_entries_barrier_2_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_2_io_y_sw = dcache_tlb_entries_barrier_2_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_sx = dcache_tlb_entries_barrier_2_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_2_io_y_sr = dcache_tlb_entries_barrier_2_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_2_io_y_hw = dcache_tlb_entries_barrier_2_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_hx = dcache_tlb_entries_barrier_2_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_2_io_y_hr = dcache_tlb_entries_barrier_2_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pw = dcache_tlb_entries_barrier_2_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_px = dcache_tlb_entries_barrier_2_io_x_px ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pr = dcache_tlb_entries_barrier_2_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ppp = dcache_tlb_entries_barrier_2_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pal = dcache_tlb_entries_barrier_2_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_2_io_y_paa = dcache_tlb_entries_barrier_2_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_2_io_y_eff = dcache_tlb_entries_barrier_2_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_2_io_y_c = dcache_tlb_entries_barrier_2_io_x_c ;
    assign  dcache_tlb_entries_barrier_3_io_y_u = dcache_tlb_entries_barrier_3_io_x_u ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ae_ptw = dcache_tlb_entries_barrier_3_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ae_final = dcache_tlb_entries_barrier_3_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ae_stage2 = dcache_tlb_entries_barrier_3_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pf = dcache_tlb_entries_barrier_3_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_3_io_y_gf = dcache_tlb_entries_barrier_3_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_3_io_y_sw = dcache_tlb_entries_barrier_3_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_sx = dcache_tlb_entries_barrier_3_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_3_io_y_sr = dcache_tlb_entries_barrier_3_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_3_io_y_hw = dcache_tlb_entries_barrier_3_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_hx = dcache_tlb_entries_barrier_3_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_3_io_y_hr = dcache_tlb_entries_barrier_3_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pw = dcache_tlb_entries_barrier_3_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_px = dcache_tlb_entries_barrier_3_io_x_px ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pr = dcache_tlb_entries_barrier_3_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ppp = dcache_tlb_entries_barrier_3_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pal = dcache_tlb_entries_barrier_3_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_3_io_y_paa = dcache_tlb_entries_barrier_3_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_3_io_y_eff = dcache_tlb_entries_barrier_3_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_3_io_y_c = dcache_tlb_entries_barrier_3_io_x_c ;
    assign  dcache_tlb_entries_barrier_4_io_y_u = dcache_tlb_entries_barrier_4_io_x_u ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ae_ptw = dcache_tlb_entries_barrier_4_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ae_final = dcache_tlb_entries_barrier_4_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ae_stage2 = dcache_tlb_entries_barrier_4_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pf = dcache_tlb_entries_barrier_4_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_4_io_y_gf = dcache_tlb_entries_barrier_4_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_4_io_y_sw = dcache_tlb_entries_barrier_4_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_sx = dcache_tlb_entries_barrier_4_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_4_io_y_sr = dcache_tlb_entries_barrier_4_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_4_io_y_hw = dcache_tlb_entries_barrier_4_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_hx = dcache_tlb_entries_barrier_4_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_4_io_y_hr = dcache_tlb_entries_barrier_4_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pw = dcache_tlb_entries_barrier_4_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_px = dcache_tlb_entries_barrier_4_io_x_px ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pr = dcache_tlb_entries_barrier_4_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ppp = dcache_tlb_entries_barrier_4_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pal = dcache_tlb_entries_barrier_4_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_4_io_y_paa = dcache_tlb_entries_barrier_4_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_4_io_y_eff = dcache_tlb_entries_barrier_4_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_4_io_y_c = dcache_tlb_entries_barrier_4_io_x_c ;
    assign  dcache_tlb_entries_barrier_5_io_y_u = dcache_tlb_entries_barrier_5_io_x_u ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ae_ptw = dcache_tlb_entries_barrier_5_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ae_final = dcache_tlb_entries_barrier_5_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ae_stage2 = dcache_tlb_entries_barrier_5_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pf = dcache_tlb_entries_barrier_5_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_5_io_y_gf = dcache_tlb_entries_barrier_5_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_5_io_y_sw = dcache_tlb_entries_barrier_5_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_sx = dcache_tlb_entries_barrier_5_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_5_io_y_sr = dcache_tlb_entries_barrier_5_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_5_io_y_hw = dcache_tlb_entries_barrier_5_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_hx = dcache_tlb_entries_barrier_5_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_5_io_y_hr = dcache_tlb_entries_barrier_5_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pw = dcache_tlb_entries_barrier_5_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_px = dcache_tlb_entries_barrier_5_io_x_px ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pr = dcache_tlb_entries_barrier_5_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ppp = dcache_tlb_entries_barrier_5_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pal = dcache_tlb_entries_barrier_5_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_5_io_y_paa = dcache_tlb_entries_barrier_5_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_5_io_y_eff = dcache_tlb_entries_barrier_5_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_5_io_y_c = dcache_tlb_entries_barrier_5_io_x_c ;
      
    
    wire dcache_pma_checker_pmp_res_cur_cfg_l = dcache_pma_checker_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_cfg_a = dcache_pma_checker_pmp_io_pmp_7_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_addr = dcache_pma_checker_pmp_io_pmp_7_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_mask = dcache_pma_checker_pmp_io_pmp_7_mask ; 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_l = dcache_pma_checker_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_1_cfg_a = dcache_pma_checker_pmp_io_pmp_6_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_1_addr = dcache_pma_checker_pmp_io_pmp_6_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_1_mask = dcache_pma_checker_pmp_io_pmp_6_mask ; 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_l = dcache_pma_checker_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_2_cfg_a = dcache_pma_checker_pmp_io_pmp_5_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_2_addr = dcache_pma_checker_pmp_io_pmp_5_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_2_mask = dcache_pma_checker_pmp_io_pmp_5_mask ; 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_l = dcache_pma_checker_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_3_cfg_a = dcache_pma_checker_pmp_io_pmp_4_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_3_addr = dcache_pma_checker_pmp_io_pmp_4_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_3_mask = dcache_pma_checker_pmp_io_pmp_4_mask ; 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_l = dcache_pma_checker_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_4_cfg_a = dcache_pma_checker_pmp_io_pmp_3_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_4_addr = dcache_pma_checker_pmp_io_pmp_3_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_4_mask = dcache_pma_checker_pmp_io_pmp_3_mask ; 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_l = dcache_pma_checker_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_5_cfg_a = dcache_pma_checker_pmp_io_pmp_2_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_5_addr = dcache_pma_checker_pmp_io_pmp_2_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_5_mask = dcache_pma_checker_pmp_io_pmp_2_mask ; 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_l = dcache_pma_checker_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_6_cfg_a = dcache_pma_checker_pmp_io_pmp_1_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_6_addr = dcache_pma_checker_pmp_io_pmp_1_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_6_mask = dcache_pma_checker_pmp_io_pmp_1_mask ; 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_l = dcache_pma_checker_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_7_cfg_a = dcache_pma_checker_pmp_io_pmp_0_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_7_addr = dcache_pma_checker_pmp_io_pmp_0_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_7_mask = dcache_pma_checker_pmp_io_pmp_0_mask ; 
    wire[1:0] dcache_pma_checker_pmp_pmp0_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_pmp0_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_1_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_2_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_3_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_4_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_5_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_6_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_7_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp_res_cfg_res =2'h0; 
    wire dcache_pma_checker_pmp_pmp0_cfg_l =1'h0; 
    wire[29:0] dcache_pma_checker_pmp_pmp0_addr =30'h0; 
    wire[31:0] dcache_pma_checker_pmp_pmp0_mask =32'h0; 
    wire dcache_pma_checker_pmp_default_0 = dcache_pma_checker_pmp_io_prv [1]; 
    wire dcache_pma_checker_pmp_pmp0_cfg_x = dcache_pma_checker_pmp_default_0 ; 
    wire dcache_pma_checker_pmp_pmp0_cfg_w = dcache_pma_checker_pmp_default_0 ; 
    wire dcache_pma_checker_pmp_pmp0_cfg_r = dcache_pma_checker_pmp_default_0 ; 
    wire dcache_pma_checker_pmp_res_hit = dcache_pma_checker_pmp_io_pmp_7_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_7_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_7_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi ; 
  assign  dcache_pma_checker_pmp_res_hi = dcache_pma_checker_pmp__GEN ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_1 ; 
  assign  dcache_pma_checker_pmp_res_hi_1 = dcache_pma_checker_pmp__GEN ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_2 ; 
  assign  dcache_pma_checker_pmp_res_hi_2 = dcache_pma_checker_pmp__GEN ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_3 ; 
  assign  dcache_pma_checker_pmp_res_hi_3 = dcache_pma_checker_pmp__GEN ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_4 ; 
  assign  dcache_pma_checker_pmp_res_hi_4 = dcache_pma_checker_pmp__GEN ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_5 ; 
  assign  dcache_pma_checker_pmp_res_hi_5 = dcache_pma_checker_pmp__GEN ; 
    wire dcache_pma_checker_pmp_res_cur_cfg_r = dcache_pma_checker_pmp_io_pmp_7_cfg_r | dcache_pma_checker_pmp_res_ignore ; 
    wire dcache_pma_checker_pmp_res_cur_cfg_w = dcache_pma_checker_pmp_io_pmp_7_cfg_w | dcache_pma_checker_pmp_res_ignore ; 
    wire dcache_pma_checker_pmp_res_cur_cfg_x = dcache_pma_checker_pmp_io_pmp_7_cfg_x | dcache_pma_checker_pmp_res_ignore ; 
    wire dcache_pma_checker_pmp_res_hit_1 = dcache_pma_checker_pmp_io_pmp_6_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_6_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_6_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_1 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_0 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_6 ; 
  assign  dcache_pma_checker_pmp_res_hi_6 = dcache_pma_checker_pmp__GEN_0 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_7 ; 
  assign  dcache_pma_checker_pmp_res_hi_7 = dcache_pma_checker_pmp__GEN_0 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_8 ; 
  assign  dcache_pma_checker_pmp_res_hi_8 = dcache_pma_checker_pmp__GEN_0 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_9 ; 
  assign  dcache_pma_checker_pmp_res_hi_9 = dcache_pma_checker_pmp__GEN_0 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_10 ; 
  assign  dcache_pma_checker_pmp_res_hi_10 = dcache_pma_checker_pmp__GEN_0 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_11 ; 
  assign  dcache_pma_checker_pmp_res_hi_11 = dcache_pma_checker_pmp__GEN_0 ; 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_r = dcache_pma_checker_pmp_io_pmp_6_cfg_r | dcache_pma_checker_pmp_res_ignore_1 ; 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_w = dcache_pma_checker_pmp_io_pmp_6_cfg_w | dcache_pma_checker_pmp_res_ignore_1 ; 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_x = dcache_pma_checker_pmp_io_pmp_6_cfg_x | dcache_pma_checker_pmp_res_ignore_1 ; 
    wire dcache_pma_checker_pmp_res_hit_2 = dcache_pma_checker_pmp_io_pmp_5_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_5_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_5_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_2 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_1 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_12 ; 
  assign  dcache_pma_checker_pmp_res_hi_12 = dcache_pma_checker_pmp__GEN_1 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_13 ; 
  assign  dcache_pma_checker_pmp_res_hi_13 = dcache_pma_checker_pmp__GEN_1 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_14 ; 
  assign  dcache_pma_checker_pmp_res_hi_14 = dcache_pma_checker_pmp__GEN_1 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_15 ; 
  assign  dcache_pma_checker_pmp_res_hi_15 = dcache_pma_checker_pmp__GEN_1 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_16 ; 
  assign  dcache_pma_checker_pmp_res_hi_16 = dcache_pma_checker_pmp__GEN_1 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_17 ; 
  assign  dcache_pma_checker_pmp_res_hi_17 = dcache_pma_checker_pmp__GEN_1 ; 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_r = dcache_pma_checker_pmp_io_pmp_5_cfg_r | dcache_pma_checker_pmp_res_ignore_2 ; 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_w = dcache_pma_checker_pmp_io_pmp_5_cfg_w | dcache_pma_checker_pmp_res_ignore_2 ; 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_x = dcache_pma_checker_pmp_io_pmp_5_cfg_x | dcache_pma_checker_pmp_res_ignore_2 ; 
    wire dcache_pma_checker_pmp_res_hit_3 = dcache_pma_checker_pmp_io_pmp_4_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_4_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_4_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_3 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_2 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_18 ; 
  assign  dcache_pma_checker_pmp_res_hi_18 = dcache_pma_checker_pmp__GEN_2 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_19 ; 
  assign  dcache_pma_checker_pmp_res_hi_19 = dcache_pma_checker_pmp__GEN_2 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_20 ; 
  assign  dcache_pma_checker_pmp_res_hi_20 = dcache_pma_checker_pmp__GEN_2 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_21 ; 
  assign  dcache_pma_checker_pmp_res_hi_21 = dcache_pma_checker_pmp__GEN_2 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_22 ; 
  assign  dcache_pma_checker_pmp_res_hi_22 = dcache_pma_checker_pmp__GEN_2 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_23 ; 
  assign  dcache_pma_checker_pmp_res_hi_23 = dcache_pma_checker_pmp__GEN_2 ; 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_r = dcache_pma_checker_pmp_io_pmp_4_cfg_r | dcache_pma_checker_pmp_res_ignore_3 ; 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_w = dcache_pma_checker_pmp_io_pmp_4_cfg_w | dcache_pma_checker_pmp_res_ignore_3 ; 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_x = dcache_pma_checker_pmp_io_pmp_4_cfg_x | dcache_pma_checker_pmp_res_ignore_3 ; 
    wire dcache_pma_checker_pmp_res_hit_4 = dcache_pma_checker_pmp_io_pmp_3_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_3_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_3_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_4 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_3 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_24 ; 
  assign  dcache_pma_checker_pmp_res_hi_24 = dcache_pma_checker_pmp__GEN_3 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_25 ; 
  assign  dcache_pma_checker_pmp_res_hi_25 = dcache_pma_checker_pmp__GEN_3 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_26 ; 
  assign  dcache_pma_checker_pmp_res_hi_26 = dcache_pma_checker_pmp__GEN_3 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_27 ; 
  assign  dcache_pma_checker_pmp_res_hi_27 = dcache_pma_checker_pmp__GEN_3 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_28 ; 
  assign  dcache_pma_checker_pmp_res_hi_28 = dcache_pma_checker_pmp__GEN_3 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_29 ; 
  assign  dcache_pma_checker_pmp_res_hi_29 = dcache_pma_checker_pmp__GEN_3 ; 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_r = dcache_pma_checker_pmp_io_pmp_3_cfg_r | dcache_pma_checker_pmp_res_ignore_4 ; 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_w = dcache_pma_checker_pmp_io_pmp_3_cfg_w | dcache_pma_checker_pmp_res_ignore_4 ; 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_x = dcache_pma_checker_pmp_io_pmp_3_cfg_x | dcache_pma_checker_pmp_res_ignore_4 ; 
    wire dcache_pma_checker_pmp_res_hit_5 = dcache_pma_checker_pmp_io_pmp_2_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_2_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_2_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_5 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_4 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_30 ; 
  assign  dcache_pma_checker_pmp_res_hi_30 = dcache_pma_checker_pmp__GEN_4 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_31 ; 
  assign  dcache_pma_checker_pmp_res_hi_31 = dcache_pma_checker_pmp__GEN_4 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_32 ; 
  assign  dcache_pma_checker_pmp_res_hi_32 = dcache_pma_checker_pmp__GEN_4 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_33 ; 
  assign  dcache_pma_checker_pmp_res_hi_33 = dcache_pma_checker_pmp__GEN_4 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_34 ; 
  assign  dcache_pma_checker_pmp_res_hi_34 = dcache_pma_checker_pmp__GEN_4 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_35 ; 
  assign  dcache_pma_checker_pmp_res_hi_35 = dcache_pma_checker_pmp__GEN_4 ; 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_r = dcache_pma_checker_pmp_io_pmp_2_cfg_r | dcache_pma_checker_pmp_res_ignore_5 ; 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_w = dcache_pma_checker_pmp_io_pmp_2_cfg_w | dcache_pma_checker_pmp_res_ignore_5 ; 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_x = dcache_pma_checker_pmp_io_pmp_2_cfg_x | dcache_pma_checker_pmp_res_ignore_5 ; 
    wire dcache_pma_checker_pmp_res_hit_6 = dcache_pma_checker_pmp_io_pmp_1_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_1_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_1_cfg_a [0]& dcache_pma_checker_pmp_io_addr >={ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_6 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_5 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_36 ; 
  assign  dcache_pma_checker_pmp_res_hi_36 = dcache_pma_checker_pmp__GEN_5 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_37 ; 
  assign  dcache_pma_checker_pmp_res_hi_37 = dcache_pma_checker_pmp__GEN_5 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_38 ; 
  assign  dcache_pma_checker_pmp_res_hi_38 = dcache_pma_checker_pmp__GEN_5 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_39 ; 
  assign  dcache_pma_checker_pmp_res_hi_39 = dcache_pma_checker_pmp__GEN_5 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_40 ; 
  assign  dcache_pma_checker_pmp_res_hi_40 = dcache_pma_checker_pmp__GEN_5 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_41 ; 
  assign  dcache_pma_checker_pmp_res_hi_41 = dcache_pma_checker_pmp__GEN_5 ; 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_r = dcache_pma_checker_pmp_io_pmp_1_cfg_r | dcache_pma_checker_pmp_res_ignore_6 ; 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_w = dcache_pma_checker_pmp_io_pmp_1_cfg_w | dcache_pma_checker_pmp_res_ignore_6 ; 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_x = dcache_pma_checker_pmp_io_pmp_1_cfg_x | dcache_pma_checker_pmp_res_ignore_6 ; 
    wire dcache_pma_checker_pmp_res_hit_7 = dcache_pma_checker_pmp_io_pmp_0_cfg_a [1] ? (( dcache_pma_checker_pmp_io_addr ^{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0})&~ dcache_pma_checker_pmp_io_pmp_0_mask )==32'h0: dcache_pma_checker_pmp_io_pmp_0_cfg_a [0]& dcache_pma_checker_pmp_io_addr <{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}; 
    wire dcache_pma_checker_pmp_res_ignore_7 = dcache_pma_checker_pmp_default_0 &~ dcache_pma_checker_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp__GEN_6 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_42 ; 
  assign  dcache_pma_checker_pmp_res_hi_42 = dcache_pma_checker_pmp__GEN_6 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_43 ; 
  assign  dcache_pma_checker_pmp_res_hi_43 = dcache_pma_checker_pmp__GEN_6 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_44 ; 
  assign  dcache_pma_checker_pmp_res_hi_44 = dcache_pma_checker_pmp__GEN_6 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_45 ; 
  assign  dcache_pma_checker_pmp_res_hi_45 = dcache_pma_checker_pmp__GEN_6 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_46 ; 
  assign  dcache_pma_checker_pmp_res_hi_46 = dcache_pma_checker_pmp__GEN_6 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_47 ; 
  assign  dcache_pma_checker_pmp_res_hi_47 = dcache_pma_checker_pmp__GEN_6 ; 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_r = dcache_pma_checker_pmp_io_pmp_0_cfg_r | dcache_pma_checker_pmp_res_ignore_7 ; 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_w = dcache_pma_checker_pmp_io_pmp_0_cfg_w | dcache_pma_checker_pmp_res_ignore_7 ; 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_x = dcache_pma_checker_pmp_io_pmp_0_cfg_x | dcache_pma_checker_pmp_res_ignore_7 ; 
    wire dcache_pma_checker_pmp_res_cfg_l = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_l : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_l : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_l : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_l : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_l : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_l : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_l : dcache_pma_checker_pmp_res_hit & dcache_pma_checker_pmp_res_cur_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cfg_a = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_a : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_a : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_a : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_a : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_a : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_a : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_a : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_a :2'h0; 
    wire dcache_pma_checker_pmp_res_cfg_x = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_x : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_x : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_x : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_x : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_x : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_x : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_x : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_x : dcache_pma_checker_pmp_pmp0_cfg_x ; 
    wire dcache_pma_checker_pmp_res_cfg_w = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_w : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_w : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_w : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_w : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_w : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_w : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_w : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_w : dcache_pma_checker_pmp_pmp0_cfg_w ; 
    wire dcache_pma_checker_pmp_res_cfg_r = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_r : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_r : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_r : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_r : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_r : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_r : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_r : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_r : dcache_pma_checker_pmp_pmp0_cfg_r ; 
    wire[29:0] dcache_pma_checker_pmp_res_addr = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_addr : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_addr : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_addr : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_addr : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_addr : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_addr : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_addr : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_addr :30'h0; 
    wire[31:0] dcache_pma_checker_pmp_res_mask = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_mask : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_mask : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_mask : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_mask : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_mask : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_mask : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_mask : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_mask :32'h0; 
  assign  dcache_pma_checker_pmp_io_r = dcache_pma_checker_pmp_res_cfg_r ; 
  assign  dcache_pma_checker_pmp_io_w = dcache_pma_checker_pmp_res_cfg_w ; 
  assign  dcache_pma_checker_pmp_io_x = dcache_pma_checker_pmp_res_cfg_x ;
    assign dcache_tlb_pmp_io_prv = dcache_tlb_mpu_priv[1:0];
    assign dcache_tlb_pmp_io_pmp_0_cfg_l = dcache_io_ptw_pmp_0_cfg_l;
    assign dcache_tlb_pmp_io_pmp_0_cfg_a = dcache_io_ptw_pmp_0_cfg_a;
    assign dcache_tlb_pmp_io_pmp_0_cfg_x = dcache_io_ptw_pmp_0_cfg_x;
    assign dcache_tlb_pmp_io_pmp_0_cfg_w = dcache_io_ptw_pmp_0_cfg_w;
    assign dcache_tlb_pmp_io_pmp_0_cfg_r = dcache_io_ptw_pmp_0_cfg_r;
    assign dcache_tlb_pmp_io_pmp_0_addr = dcache_io_ptw_pmp_0_addr;
    assign dcache_tlb_pmp_io_pmp_0_mask = dcache_io_ptw_pmp_0_mask;
    assign dcache_tlb_pmp_io_pmp_1_cfg_l = dcache_io_ptw_pmp_1_cfg_l;
    assign dcache_tlb_pmp_io_pmp_1_cfg_a = dcache_io_ptw_pmp_1_cfg_a;
    assign dcache_tlb_pmp_io_pmp_1_cfg_x = dcache_io_ptw_pmp_1_cfg_x;
    assign dcache_tlb_pmp_io_pmp_1_cfg_w = dcache_io_ptw_pmp_1_cfg_w;
    assign dcache_tlb_pmp_io_pmp_1_cfg_r = dcache_io_ptw_pmp_1_cfg_r;
    assign dcache_tlb_pmp_io_pmp_1_addr = dcache_io_ptw_pmp_1_addr;
    assign dcache_tlb_pmp_io_pmp_1_mask = dcache_io_ptw_pmp_1_mask;
    assign dcache_tlb_pmp_io_pmp_2_cfg_l = dcache_io_ptw_pmp_2_cfg_l;
    assign dcache_tlb_pmp_io_pmp_2_cfg_a = dcache_io_ptw_pmp_2_cfg_a;
    assign dcache_tlb_pmp_io_pmp_2_cfg_x = dcache_io_ptw_pmp_2_cfg_x;
    assign dcache_tlb_pmp_io_pmp_2_cfg_w = dcache_io_ptw_pmp_2_cfg_w;
    assign dcache_tlb_pmp_io_pmp_2_cfg_r = dcache_io_ptw_pmp_2_cfg_r;
    assign dcache_tlb_pmp_io_pmp_2_addr = dcache_io_ptw_pmp_2_addr;
    assign dcache_tlb_pmp_io_pmp_2_mask = dcache_io_ptw_pmp_2_mask;
    assign dcache_tlb_pmp_io_pmp_3_cfg_l = dcache_io_ptw_pmp_3_cfg_l;
    assign dcache_tlb_pmp_io_pmp_3_cfg_a = dcache_io_ptw_pmp_3_cfg_a;
    assign dcache_tlb_pmp_io_pmp_3_cfg_x = dcache_io_ptw_pmp_3_cfg_x;
    assign dcache_tlb_pmp_io_pmp_3_cfg_w = dcache_io_ptw_pmp_3_cfg_w;
    assign dcache_tlb_pmp_io_pmp_3_cfg_r = dcache_io_ptw_pmp_3_cfg_r;
    assign dcache_tlb_pmp_io_pmp_3_addr = dcache_io_ptw_pmp_3_addr;
    assign dcache_tlb_pmp_io_pmp_3_mask = dcache_io_ptw_pmp_3_mask;
    assign dcache_tlb_pmp_io_pmp_4_cfg_l = dcache_io_ptw_pmp_4_cfg_l;
    assign dcache_tlb_pmp_io_pmp_4_cfg_a = dcache_io_ptw_pmp_4_cfg_a;
    assign dcache_tlb_pmp_io_pmp_4_cfg_x = dcache_io_ptw_pmp_4_cfg_x;
    assign dcache_tlb_pmp_io_pmp_4_cfg_w = dcache_io_ptw_pmp_4_cfg_w;
    assign dcache_tlb_pmp_io_pmp_4_cfg_r = dcache_io_ptw_pmp_4_cfg_r;
    assign dcache_tlb_pmp_io_pmp_4_addr = dcache_io_ptw_pmp_4_addr;
    assign dcache_tlb_pmp_io_pmp_4_mask = dcache_io_ptw_pmp_4_mask;
    assign dcache_tlb_pmp_io_pmp_5_cfg_l = dcache_io_ptw_pmp_5_cfg_l;
    assign dcache_tlb_pmp_io_pmp_5_cfg_a = dcache_io_ptw_pmp_5_cfg_a;
    assign dcache_tlb_pmp_io_pmp_5_cfg_x = dcache_io_ptw_pmp_5_cfg_x;
    assign dcache_tlb_pmp_io_pmp_5_cfg_w = dcache_io_ptw_pmp_5_cfg_w;
    assign dcache_tlb_pmp_io_pmp_5_cfg_r = dcache_io_ptw_pmp_5_cfg_r;
    assign dcache_tlb_pmp_io_pmp_5_addr = dcache_io_ptw_pmp_5_addr;
    assign dcache_tlb_pmp_io_pmp_5_mask = dcache_io_ptw_pmp_5_mask;
    assign dcache_tlb_pmp_io_pmp_6_cfg_l = dcache_io_ptw_pmp_6_cfg_l;
    assign dcache_tlb_pmp_io_pmp_6_cfg_a = dcache_io_ptw_pmp_6_cfg_a;
    assign dcache_tlb_pmp_io_pmp_6_cfg_x = dcache_io_ptw_pmp_6_cfg_x;
    assign dcache_tlb_pmp_io_pmp_6_cfg_w = dcache_io_ptw_pmp_6_cfg_w;
    assign dcache_tlb_pmp_io_pmp_6_cfg_r = dcache_io_ptw_pmp_6_cfg_r;
    assign dcache_tlb_pmp_io_pmp_6_addr = dcache_io_ptw_pmp_6_addr;
    assign dcache_tlb_pmp_io_pmp_6_mask = dcache_io_ptw_pmp_6_mask;
    assign dcache_tlb_pmp_io_pmp_7_cfg_l = dcache_io_ptw_pmp_7_cfg_l;
    assign dcache_tlb_pmp_io_pmp_7_cfg_a = dcache_io_ptw_pmp_7_cfg_a;
    assign dcache_tlb_pmp_io_pmp_7_cfg_x = dcache_io_ptw_pmp_7_cfg_x;
    assign dcache_tlb_pmp_io_pmp_7_cfg_w = dcache_io_ptw_pmp_7_cfg_w;
    assign dcache_tlb_pmp_io_pmp_7_cfg_r = dcache_io_ptw_pmp_7_cfg_r;
    assign dcache_tlb_pmp_io_pmp_7_addr = dcache_io_ptw_pmp_7_addr;
    assign dcache_tlb_pmp_io_pmp_7_mask = dcache_io_ptw_pmp_7_mask;
    assign dcache_tlb_pmp_io_addr = dcache_tlb_mpu_physaddr;
    assign dcache__tlb_pmp_io_r = dcache_tlb_pmp_io_r;
    assign dcache__tlb_pmp_io_w = dcache_tlb_pmp_io_w;
    assign dcache__tlb_pmp_io_x = dcache_tlb_pmp_io_x;
    assign dcache_pma_checker_pmp_io_prv = dcache_pma_checker_mpu_priv[1:0];
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_0_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_0_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_1_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_2_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_3_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_4_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_5_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_6_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_l = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_a = 2'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_x = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_w = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_r = 1'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_addr = 30'h0;
    assign dcache_pma_checker_pmp_io_pmp_7_mask = 32'h0;
    assign dcache_pma_checker_pmp_io_addr = dcache_pma_checker_mpu_physaddr;
    assign dcache__pma_checker_pmp_io_r = dcache_pma_checker_pmp_io_r;
    assign dcache__pma_checker_pmp_io_w = dcache_pma_checker_pmp_io_w;
    assign dcache__pma_checker_pmp_io_x = dcache_pma_checker_pmp_io_x;
      
    
    assign  dcache_pma_checker_entries_barrier_io_y_u = dcache_pma_checker_entries_barrier_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ae_ptw = dcache_pma_checker_entries_barrier_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ae_final = dcache_pma_checker_entries_barrier_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pf = dcache_pma_checker_entries_barrier_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_io_y_gf = dcache_pma_checker_entries_barrier_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_io_y_sw = dcache_pma_checker_entries_barrier_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_sx = dcache_pma_checker_entries_barrier_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_io_y_sr = dcache_pma_checker_entries_barrier_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_io_y_hw = dcache_pma_checker_entries_barrier_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_hx = dcache_pma_checker_entries_barrier_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_io_y_hr = dcache_pma_checker_entries_barrier_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pw = dcache_pma_checker_entries_barrier_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_px = dcache_pma_checker_entries_barrier_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pr = dcache_pma_checker_entries_barrier_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ppp = dcache_pma_checker_entries_barrier_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pal = dcache_pma_checker_entries_barrier_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_io_y_paa = dcache_pma_checker_entries_barrier_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_io_y_eff = dcache_pma_checker_entries_barrier_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_io_y_c = dcache_pma_checker_entries_barrier_io_x_c ;
    assign  dcache_pma_checker_entries_barrier_1_io_y_u = dcache_pma_checker_entries_barrier_1_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ae_ptw = dcache_pma_checker_entries_barrier_1_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ae_final = dcache_pma_checker_entries_barrier_1_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_1_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pf = dcache_pma_checker_entries_barrier_1_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_gf = dcache_pma_checker_entries_barrier_1_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_sw = dcache_pma_checker_entries_barrier_1_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_sx = dcache_pma_checker_entries_barrier_1_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_sr = dcache_pma_checker_entries_barrier_1_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_hw = dcache_pma_checker_entries_barrier_1_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_hx = dcache_pma_checker_entries_barrier_1_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_hr = dcache_pma_checker_entries_barrier_1_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pw = dcache_pma_checker_entries_barrier_1_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_px = dcache_pma_checker_entries_barrier_1_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pr = dcache_pma_checker_entries_barrier_1_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ppp = dcache_pma_checker_entries_barrier_1_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pal = dcache_pma_checker_entries_barrier_1_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_paa = dcache_pma_checker_entries_barrier_1_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_eff = dcache_pma_checker_entries_barrier_1_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_c = dcache_pma_checker_entries_barrier_1_io_x_c ;
    assign  dcache_pma_checker_entries_barrier_2_io_y_u = dcache_pma_checker_entries_barrier_2_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ae_ptw = dcache_pma_checker_entries_barrier_2_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ae_final = dcache_pma_checker_entries_barrier_2_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_2_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pf = dcache_pma_checker_entries_barrier_2_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_gf = dcache_pma_checker_entries_barrier_2_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_sw = dcache_pma_checker_entries_barrier_2_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_sx = dcache_pma_checker_entries_barrier_2_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_sr = dcache_pma_checker_entries_barrier_2_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_hw = dcache_pma_checker_entries_barrier_2_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_hx = dcache_pma_checker_entries_barrier_2_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_hr = dcache_pma_checker_entries_barrier_2_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pw = dcache_pma_checker_entries_barrier_2_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_px = dcache_pma_checker_entries_barrier_2_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pr = dcache_pma_checker_entries_barrier_2_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ppp = dcache_pma_checker_entries_barrier_2_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pal = dcache_pma_checker_entries_barrier_2_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_paa = dcache_pma_checker_entries_barrier_2_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_eff = dcache_pma_checker_entries_barrier_2_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_c = dcache_pma_checker_entries_barrier_2_io_x_c ;
    assign  dcache_pma_checker_entries_barrier_3_io_y_u = dcache_pma_checker_entries_barrier_3_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ae_ptw = dcache_pma_checker_entries_barrier_3_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ae_final = dcache_pma_checker_entries_barrier_3_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_3_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pf = dcache_pma_checker_entries_barrier_3_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_gf = dcache_pma_checker_entries_barrier_3_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_sw = dcache_pma_checker_entries_barrier_3_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_sx = dcache_pma_checker_entries_barrier_3_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_sr = dcache_pma_checker_entries_barrier_3_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_hw = dcache_pma_checker_entries_barrier_3_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_hx = dcache_pma_checker_entries_barrier_3_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_hr = dcache_pma_checker_entries_barrier_3_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pw = dcache_pma_checker_entries_barrier_3_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_px = dcache_pma_checker_entries_barrier_3_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pr = dcache_pma_checker_entries_barrier_3_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ppp = dcache_pma_checker_entries_barrier_3_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pal = dcache_pma_checker_entries_barrier_3_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_paa = dcache_pma_checker_entries_barrier_3_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_eff = dcache_pma_checker_entries_barrier_3_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_c = dcache_pma_checker_entries_barrier_3_io_x_c ;
    assign  dcache_pma_checker_entries_barrier_4_io_y_u = dcache_pma_checker_entries_barrier_4_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ae_ptw = dcache_pma_checker_entries_barrier_4_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ae_final = dcache_pma_checker_entries_barrier_4_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_4_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pf = dcache_pma_checker_entries_barrier_4_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_gf = dcache_pma_checker_entries_barrier_4_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_sw = dcache_pma_checker_entries_barrier_4_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_sx = dcache_pma_checker_entries_barrier_4_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_sr = dcache_pma_checker_entries_barrier_4_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_hw = dcache_pma_checker_entries_barrier_4_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_hx = dcache_pma_checker_entries_barrier_4_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_hr = dcache_pma_checker_entries_barrier_4_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pw = dcache_pma_checker_entries_barrier_4_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_px = dcache_pma_checker_entries_barrier_4_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pr = dcache_pma_checker_entries_barrier_4_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ppp = dcache_pma_checker_entries_barrier_4_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pal = dcache_pma_checker_entries_barrier_4_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_paa = dcache_pma_checker_entries_barrier_4_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_eff = dcache_pma_checker_entries_barrier_4_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_c = dcache_pma_checker_entries_barrier_4_io_x_c ;
    assign  dcache_pma_checker_entries_barrier_5_io_y_u = dcache_pma_checker_entries_barrier_5_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ae_ptw = dcache_pma_checker_entries_barrier_5_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ae_final = dcache_pma_checker_entries_barrier_5_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_5_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pf = dcache_pma_checker_entries_barrier_5_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_gf = dcache_pma_checker_entries_barrier_5_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_sw = dcache_pma_checker_entries_barrier_5_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_sx = dcache_pma_checker_entries_barrier_5_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_sr = dcache_pma_checker_entries_barrier_5_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_hw = dcache_pma_checker_entries_barrier_5_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_hx = dcache_pma_checker_entries_barrier_5_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_hr = dcache_pma_checker_entries_barrier_5_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pw = dcache_pma_checker_entries_barrier_5_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_px = dcache_pma_checker_entries_barrier_5_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pr = dcache_pma_checker_entries_barrier_5_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ppp = dcache_pma_checker_entries_barrier_5_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pal = dcache_pma_checker_entries_barrier_5_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_paa = dcache_pma_checker_entries_barrier_5_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_eff = dcache_pma_checker_entries_barrier_5_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_c = dcache_pma_checker_entries_barrier_5_io_x_c ;
    assign dcache_tlb_entries_barrier_io_x_u = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_ae_ptw = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_ae_final = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_ae_stage2 = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_pf = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_gf = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_sw = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_sx = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_sr = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_hw = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_hx = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_hr = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_pw = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_px = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_pr = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_ppp = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_pal = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_paa = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_eff = 1'h0;
    assign dcache_tlb_entries_barrier_io_x_c = 1'h0;
    assign dcache__tlb_entries_barrier_io_y_u = dcache_tlb_entries_barrier_io_y_u;
    assign dcache__tlb_entries_barrier_io_y_ae_ptw = dcache_tlb_entries_barrier_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_io_y_ae_final = dcache_tlb_entries_barrier_io_y_ae_final;
    assign dcache__tlb_entries_barrier_io_y_ae_stage2 = dcache_tlb_entries_barrier_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_io_y_pf = dcache_tlb_entries_barrier_io_y_pf;
    assign dcache__tlb_entries_barrier_io_y_gf = dcache_tlb_entries_barrier_io_y_gf;
    assign dcache__tlb_entries_barrier_io_y_sw = dcache_tlb_entries_barrier_io_y_sw;
    assign dcache__tlb_entries_barrier_io_y_sx = dcache_tlb_entries_barrier_io_y_sx;
    assign dcache__tlb_entries_barrier_io_y_sr = dcache_tlb_entries_barrier_io_y_sr;
    assign dcache__tlb_entries_barrier_io_y_hw = dcache_tlb_entries_barrier_io_y_hw;
    assign dcache__tlb_entries_barrier_io_y_hx = dcache_tlb_entries_barrier_io_y_hx;
    assign dcache__tlb_entries_barrier_io_y_hr = dcache_tlb_entries_barrier_io_y_hr;
    assign dcache__tlb_entries_barrier_io_y_pw = dcache_tlb_entries_barrier_io_y_pw;
    assign dcache__tlb_entries_barrier_io_y_px = dcache_tlb_entries_barrier_io_y_px;
    assign dcache__tlb_entries_barrier_io_y_pr = dcache_tlb_entries_barrier_io_y_pr;
    assign dcache__tlb_entries_barrier_io_y_ppp = dcache_tlb_entries_barrier_io_y_ppp;
    assign dcache__tlb_entries_barrier_io_y_pal = dcache_tlb_entries_barrier_io_y_pal;
    assign dcache__tlb_entries_barrier_io_y_paa = dcache_tlb_entries_barrier_io_y_paa;
    assign dcache__tlb_entries_barrier_io_y_eff = dcache_tlb_entries_barrier_io_y_eff;
    assign dcache__tlb_entries_barrier_io_y_c = dcache_tlb_entries_barrier_io_y_c;
    assign dcache_tlb_entries_barrier_1_io_x_u = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_ae_ptw = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_ae_final = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_ae_stage2 = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_pf = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_gf = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_sw = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_sx = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_sr = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_hw = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_hx = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_hr = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_pw = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_px = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_pr = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_ppp = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_pal = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_paa = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_eff = 1'h0;
    assign dcache_tlb_entries_barrier_1_io_x_c = 1'h0;
    assign dcache__tlb_entries_barrier_1_io_y_u = dcache_tlb_entries_barrier_1_io_y_u;
    assign dcache__tlb_entries_barrier_1_io_y_ae_ptw = dcache_tlb_entries_barrier_1_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_1_io_y_ae_final = dcache_tlb_entries_barrier_1_io_y_ae_final;
    assign dcache__tlb_entries_barrier_1_io_y_ae_stage2 = dcache_tlb_entries_barrier_1_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_1_io_y_pf = dcache_tlb_entries_barrier_1_io_y_pf;
    assign dcache__tlb_entries_barrier_1_io_y_gf = dcache_tlb_entries_barrier_1_io_y_gf;
    assign dcache__tlb_entries_barrier_1_io_y_sw = dcache_tlb_entries_barrier_1_io_y_sw;
    assign dcache__tlb_entries_barrier_1_io_y_sx = dcache_tlb_entries_barrier_1_io_y_sx;
    assign dcache__tlb_entries_barrier_1_io_y_sr = dcache_tlb_entries_barrier_1_io_y_sr;
    assign dcache__tlb_entries_barrier_1_io_y_hw = dcache_tlb_entries_barrier_1_io_y_hw;
    assign dcache__tlb_entries_barrier_1_io_y_hx = dcache_tlb_entries_barrier_1_io_y_hx;
    assign dcache__tlb_entries_barrier_1_io_y_hr = dcache_tlb_entries_barrier_1_io_y_hr;
    assign dcache__tlb_entries_barrier_1_io_y_pw = dcache_tlb_entries_barrier_1_io_y_pw;
    assign dcache__tlb_entries_barrier_1_io_y_px = dcache_tlb_entries_barrier_1_io_y_px;
    assign dcache__tlb_entries_barrier_1_io_y_pr = dcache_tlb_entries_barrier_1_io_y_pr;
    assign dcache__tlb_entries_barrier_1_io_y_ppp = dcache_tlb_entries_barrier_1_io_y_ppp;
    assign dcache__tlb_entries_barrier_1_io_y_pal = dcache_tlb_entries_barrier_1_io_y_pal;
    assign dcache__tlb_entries_barrier_1_io_y_paa = dcache_tlb_entries_barrier_1_io_y_paa;
    assign dcache__tlb_entries_barrier_1_io_y_eff = dcache_tlb_entries_barrier_1_io_y_eff;
    assign dcache__tlb_entries_barrier_1_io_y_c = dcache_tlb_entries_barrier_1_io_y_c;
    assign dcache_tlb_entries_barrier_2_io_x_u = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_ae_ptw = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_ae_final = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_ae_stage2 = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_pf = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_gf = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_sw = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_sx = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_sr = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_hw = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_hx = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_hr = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_pw = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_px = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_pr = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_ppp = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_pal = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_paa = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_eff = 1'h0;
    assign dcache_tlb_entries_barrier_2_io_x_c = 1'h0;
    assign dcache__tlb_entries_barrier_2_io_y_u = dcache_tlb_entries_barrier_2_io_y_u;
    assign dcache__tlb_entries_barrier_2_io_y_ae_ptw = dcache_tlb_entries_barrier_2_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_2_io_y_ae_final = dcache_tlb_entries_barrier_2_io_y_ae_final;
    assign dcache__tlb_entries_barrier_2_io_y_ae_stage2 = dcache_tlb_entries_barrier_2_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_2_io_y_pf = dcache_tlb_entries_barrier_2_io_y_pf;
    assign dcache__tlb_entries_barrier_2_io_y_gf = dcache_tlb_entries_barrier_2_io_y_gf;
    assign dcache__tlb_entries_barrier_2_io_y_sw = dcache_tlb_entries_barrier_2_io_y_sw;
    assign dcache__tlb_entries_barrier_2_io_y_sx = dcache_tlb_entries_barrier_2_io_y_sx;
    assign dcache__tlb_entries_barrier_2_io_y_sr = dcache_tlb_entries_barrier_2_io_y_sr;
    assign dcache__tlb_entries_barrier_2_io_y_hw = dcache_tlb_entries_barrier_2_io_y_hw;
    assign dcache__tlb_entries_barrier_2_io_y_hx = dcache_tlb_entries_barrier_2_io_y_hx;
    assign dcache__tlb_entries_barrier_2_io_y_hr = dcache_tlb_entries_barrier_2_io_y_hr;
    assign dcache__tlb_entries_barrier_2_io_y_pw = dcache_tlb_entries_barrier_2_io_y_pw;
    assign dcache__tlb_entries_barrier_2_io_y_px = dcache_tlb_entries_barrier_2_io_y_px;
    assign dcache__tlb_entries_barrier_2_io_y_pr = dcache_tlb_entries_barrier_2_io_y_pr;
    assign dcache__tlb_entries_barrier_2_io_y_ppp = dcache_tlb_entries_barrier_2_io_y_ppp;
    assign dcache__tlb_entries_barrier_2_io_y_pal = dcache_tlb_entries_barrier_2_io_y_pal;
    assign dcache__tlb_entries_barrier_2_io_y_paa = dcache_tlb_entries_barrier_2_io_y_paa;
    assign dcache__tlb_entries_barrier_2_io_y_eff = dcache_tlb_entries_barrier_2_io_y_eff;
    assign dcache__tlb_entries_barrier_2_io_y_c = dcache_tlb_entries_barrier_2_io_y_c;
    assign dcache_tlb_entries_barrier_3_io_x_u = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_ae_ptw = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_ae_final = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_ae_stage2 = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_pf = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_gf = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_sw = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_sx = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_sr = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_hw = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_hx = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_hr = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_pw = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_px = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_pr = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_ppp = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_pal = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_paa = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_eff = 1'h0;
    assign dcache_tlb_entries_barrier_3_io_x_c = 1'h0;
    assign dcache__tlb_entries_barrier_3_io_y_u = dcache_tlb_entries_barrier_3_io_y_u;
    assign dcache__tlb_entries_barrier_3_io_y_ae_ptw = dcache_tlb_entries_barrier_3_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_3_io_y_ae_final = dcache_tlb_entries_barrier_3_io_y_ae_final;
    assign dcache__tlb_entries_barrier_3_io_y_ae_stage2 = dcache_tlb_entries_barrier_3_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_3_io_y_pf = dcache_tlb_entries_barrier_3_io_y_pf;
    assign dcache__tlb_entries_barrier_3_io_y_gf = dcache_tlb_entries_barrier_3_io_y_gf;
    assign dcache__tlb_entries_barrier_3_io_y_sw = dcache_tlb_entries_barrier_3_io_y_sw;
    assign dcache__tlb_entries_barrier_3_io_y_sx = dcache_tlb_entries_barrier_3_io_y_sx;
    assign dcache__tlb_entries_barrier_3_io_y_sr = dcache_tlb_entries_barrier_3_io_y_sr;
    assign dcache__tlb_entries_barrier_3_io_y_hw = dcache_tlb_entries_barrier_3_io_y_hw;
    assign dcache__tlb_entries_barrier_3_io_y_hx = dcache_tlb_entries_barrier_3_io_y_hx;
    assign dcache__tlb_entries_barrier_3_io_y_hr = dcache_tlb_entries_barrier_3_io_y_hr;
    assign dcache__tlb_entries_barrier_3_io_y_pw = dcache_tlb_entries_barrier_3_io_y_pw;
    assign dcache__tlb_entries_barrier_3_io_y_px = dcache_tlb_entries_barrier_3_io_y_px;
    assign dcache__tlb_entries_barrier_3_io_y_pr = dcache_tlb_entries_barrier_3_io_y_pr;
    assign dcache__tlb_entries_barrier_3_io_y_ppp = dcache_tlb_entries_barrier_3_io_y_ppp;
    assign dcache__tlb_entries_barrier_3_io_y_pal = dcache_tlb_entries_barrier_3_io_y_pal;
    assign dcache__tlb_entries_barrier_3_io_y_paa = dcache_tlb_entries_barrier_3_io_y_paa;
    assign dcache__tlb_entries_barrier_3_io_y_eff = dcache_tlb_entries_barrier_3_io_y_eff;
    assign dcache__tlb_entries_barrier_3_io_y_c = dcache_tlb_entries_barrier_3_io_y_c;
    assign dcache_tlb_entries_barrier_4_io_x_u = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_ae_ptw = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_ae_final = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_ae_stage2 = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_pf = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_gf = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_sw = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_sx = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_sr = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_hw = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_hx = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_hr = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_pw = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_px = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_pr = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_ppp = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_pal = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_paa = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_eff = 1'h0;
    assign dcache_tlb_entries_barrier_4_io_x_c = 1'h0;
    assign dcache__tlb_entries_barrier_4_io_y_u = dcache_tlb_entries_barrier_4_io_y_u;
    assign dcache__tlb_entries_barrier_4_io_y_ae_ptw = dcache_tlb_entries_barrier_4_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_4_io_y_ae_final = dcache_tlb_entries_barrier_4_io_y_ae_final;
    assign dcache__tlb_entries_barrier_4_io_y_ae_stage2 = dcache_tlb_entries_barrier_4_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_4_io_y_pf = dcache_tlb_entries_barrier_4_io_y_pf;
    assign dcache__tlb_entries_barrier_4_io_y_gf = dcache_tlb_entries_barrier_4_io_y_gf;
    assign dcache__tlb_entries_barrier_4_io_y_sw = dcache_tlb_entries_barrier_4_io_y_sw;
    assign dcache__tlb_entries_barrier_4_io_y_sx = dcache_tlb_entries_barrier_4_io_y_sx;
    assign dcache__tlb_entries_barrier_4_io_y_sr = dcache_tlb_entries_barrier_4_io_y_sr;
    assign dcache__tlb_entries_barrier_4_io_y_hw = dcache_tlb_entries_barrier_4_io_y_hw;
    assign dcache__tlb_entries_barrier_4_io_y_hx = dcache_tlb_entries_barrier_4_io_y_hx;
    assign dcache__tlb_entries_barrier_4_io_y_hr = dcache_tlb_entries_barrier_4_io_y_hr;
    assign dcache__tlb_entries_barrier_4_io_y_pw = dcache_tlb_entries_barrier_4_io_y_pw;
    assign dcache__tlb_entries_barrier_4_io_y_px = dcache_tlb_entries_barrier_4_io_y_px;
    assign dcache__tlb_entries_barrier_4_io_y_pr = dcache_tlb_entries_barrier_4_io_y_pr;
    assign dcache__tlb_entries_barrier_4_io_y_ppp = dcache_tlb_entries_barrier_4_io_y_ppp;
    assign dcache__tlb_entries_barrier_4_io_y_pal = dcache_tlb_entries_barrier_4_io_y_pal;
    assign dcache__tlb_entries_barrier_4_io_y_paa = dcache_tlb_entries_barrier_4_io_y_paa;
    assign dcache__tlb_entries_barrier_4_io_y_eff = dcache_tlb_entries_barrier_4_io_y_eff;
    assign dcache__tlb_entries_barrier_4_io_y_c = dcache_tlb_entries_barrier_4_io_y_c;
    assign dcache_tlb_entries_barrier_5_io_x_u = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_ae_ptw = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_ae_final = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_ae_stage2 = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_pf = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_gf = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_sw = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_sx = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_sr = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_hw = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_hx = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_hr = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_pw = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_px = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_pr = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_ppp = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_pal = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_paa = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_eff = 1'h0;
    assign dcache_tlb_entries_barrier_5_io_x_c = 1'h0;
    assign dcache__tlb_entries_barrier_5_io_y_u = dcache_tlb_entries_barrier_5_io_y_u;
    assign dcache__tlb_entries_barrier_5_io_y_ae_ptw = dcache_tlb_entries_barrier_5_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_5_io_y_ae_final = dcache_tlb_entries_barrier_5_io_y_ae_final;
    assign dcache__tlb_entries_barrier_5_io_y_ae_stage2 = dcache_tlb_entries_barrier_5_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_5_io_y_pf = dcache_tlb_entries_barrier_5_io_y_pf;
    assign dcache__tlb_entries_barrier_5_io_y_gf = dcache_tlb_entries_barrier_5_io_y_gf;
    assign dcache__tlb_entries_barrier_5_io_y_sw = dcache_tlb_entries_barrier_5_io_y_sw;
    assign dcache__tlb_entries_barrier_5_io_y_sx = dcache_tlb_entries_barrier_5_io_y_sx;
    assign dcache__tlb_entries_barrier_5_io_y_sr = dcache_tlb_entries_barrier_5_io_y_sr;
    assign dcache__tlb_entries_barrier_5_io_y_hw = dcache_tlb_entries_barrier_5_io_y_hw;
    assign dcache__tlb_entries_barrier_5_io_y_hx = dcache_tlb_entries_barrier_5_io_y_hx;
    assign dcache__tlb_entries_barrier_5_io_y_hr = dcache_tlb_entries_barrier_5_io_y_hr;
    assign dcache_pma_checker_entries_barrier_io_x_u = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_ae_ptw = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_ae_final = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_ae_stage2 = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_pf = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_gf = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_sw = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_sx = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_sr = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_hw = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_hx = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_hr = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_pw = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_px = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_pr = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_ppp = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_pal = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_paa = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_eff = 1'h0;
    assign dcache_pma_checker_entries_barrier_io_x_c = 1'h0;
    assign dcache__pma_checker_entries_barrier_io_y_u = dcache_pma_checker_entries_barrier_io_y_u;
    assign dcache__pma_checker_entries_barrier_io_y_ae_ptw = dcache_pma_checker_entries_barrier_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_io_y_ae_final = dcache_pma_checker_entries_barrier_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_io_y_pf = dcache_pma_checker_entries_barrier_io_y_pf;
    assign dcache__pma_checker_entries_barrier_io_y_gf = dcache_pma_checker_entries_barrier_io_y_gf;
    assign dcache__pma_checker_entries_barrier_io_y_sw = dcache_pma_checker_entries_barrier_io_y_sw;
    assign dcache__pma_checker_entries_barrier_io_y_sx = dcache_pma_checker_entries_barrier_io_y_sx;
    assign dcache__pma_checker_entries_barrier_io_y_sr = dcache_pma_checker_entries_barrier_io_y_sr;
    assign dcache__pma_checker_entries_barrier_io_y_hw = dcache_pma_checker_entries_barrier_io_y_hw;
    assign dcache__pma_checker_entries_barrier_io_y_hx = dcache_pma_checker_entries_barrier_io_y_hx;
    assign dcache__pma_checker_entries_barrier_io_y_hr = dcache_pma_checker_entries_barrier_io_y_hr;
    assign dcache__pma_checker_entries_barrier_io_y_pw = dcache_pma_checker_entries_barrier_io_y_pw;
    assign dcache__pma_checker_entries_barrier_io_y_px = dcache_pma_checker_entries_barrier_io_y_px;
    assign dcache__pma_checker_entries_barrier_io_y_pr = dcache_pma_checker_entries_barrier_io_y_pr;
    assign dcache__pma_checker_entries_barrier_io_y_ppp = dcache_pma_checker_entries_barrier_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_io_y_pal = dcache_pma_checker_entries_barrier_io_y_pal;
    assign dcache__pma_checker_entries_barrier_io_y_paa = dcache_pma_checker_entries_barrier_io_y_paa;
    assign dcache__pma_checker_entries_barrier_io_y_eff = dcache_pma_checker_entries_barrier_io_y_eff;
    assign dcache__pma_checker_entries_barrier_io_y_c = dcache_pma_checker_entries_barrier_io_y_c;
    assign dcache_pma_checker_entries_barrier_1_io_x_u = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_ae_ptw = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_ae_final = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_ae_stage2 = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_pf = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_gf = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_sw = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_sx = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_sr = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_hw = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_hx = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_hr = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_pw = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_px = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_pr = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_ppp = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_pal = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_paa = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_eff = 1'h0;
    assign dcache_pma_checker_entries_barrier_1_io_x_c = 1'h0;
    assign dcache__pma_checker_entries_barrier_1_io_y_u = dcache_pma_checker_entries_barrier_1_io_y_u;
    assign dcache__pma_checker_entries_barrier_1_io_y_ae_ptw = dcache_pma_checker_entries_barrier_1_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_1_io_y_ae_final = dcache_pma_checker_entries_barrier_1_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_1_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_1_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_1_io_y_pf = dcache_pma_checker_entries_barrier_1_io_y_pf;
    assign dcache__pma_checker_entries_barrier_1_io_y_gf = dcache_pma_checker_entries_barrier_1_io_y_gf;
    assign dcache__pma_checker_entries_barrier_1_io_y_sw = dcache_pma_checker_entries_barrier_1_io_y_sw;
    assign dcache__pma_checker_entries_barrier_1_io_y_sx = dcache_pma_checker_entries_barrier_1_io_y_sx;
    assign dcache__pma_checker_entries_barrier_1_io_y_sr = dcache_pma_checker_entries_barrier_1_io_y_sr;
    assign dcache__pma_checker_entries_barrier_1_io_y_hw = dcache_pma_checker_entries_barrier_1_io_y_hw;
    assign dcache__pma_checker_entries_barrier_1_io_y_hx = dcache_pma_checker_entries_barrier_1_io_y_hx;
    assign dcache__pma_checker_entries_barrier_1_io_y_hr = dcache_pma_checker_entries_barrier_1_io_y_hr;
    assign dcache__pma_checker_entries_barrier_1_io_y_pw = dcache_pma_checker_entries_barrier_1_io_y_pw;
    assign dcache__pma_checker_entries_barrier_1_io_y_px = dcache_pma_checker_entries_barrier_1_io_y_px;
    assign dcache__pma_checker_entries_barrier_1_io_y_pr = dcache_pma_checker_entries_barrier_1_io_y_pr;
    assign dcache__pma_checker_entries_barrier_1_io_y_ppp = dcache_pma_checker_entries_barrier_1_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_1_io_y_pal = dcache_pma_checker_entries_barrier_1_io_y_pal;
    assign dcache__pma_checker_entries_barrier_1_io_y_paa = dcache_pma_checker_entries_barrier_1_io_y_paa;
    assign dcache__pma_checker_entries_barrier_1_io_y_eff = dcache_pma_checker_entries_barrier_1_io_y_eff;
    assign dcache__pma_checker_entries_barrier_1_io_y_c = dcache_pma_checker_entries_barrier_1_io_y_c;
    assign dcache_pma_checker_entries_barrier_2_io_x_u = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_ae_ptw = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_ae_final = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_ae_stage2 = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_pf = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_gf = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_sw = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_sx = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_sr = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_hw = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_hx = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_hr = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_pw = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_px = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_pr = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_ppp = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_pal = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_paa = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_eff = 1'h0;
    assign dcache_pma_checker_entries_barrier_2_io_x_c = 1'h0;
    assign dcache__pma_checker_entries_barrier_2_io_y_u = dcache_pma_checker_entries_barrier_2_io_y_u;
    assign dcache__pma_checker_entries_barrier_2_io_y_ae_ptw = dcache_pma_checker_entries_barrier_2_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_2_io_y_ae_final = dcache_pma_checker_entries_barrier_2_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_2_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_2_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_2_io_y_pf = dcache_pma_checker_entries_barrier_2_io_y_pf;
    assign dcache__pma_checker_entries_barrier_2_io_y_gf = dcache_pma_checker_entries_barrier_2_io_y_gf;
    assign dcache__pma_checker_entries_barrier_2_io_y_sw = dcache_pma_checker_entries_barrier_2_io_y_sw;
    assign dcache__pma_checker_entries_barrier_2_io_y_sx = dcache_pma_checker_entries_barrier_2_io_y_sx;
    assign dcache__pma_checker_entries_barrier_2_io_y_sr = dcache_pma_checker_entries_barrier_2_io_y_sr;
    assign dcache__pma_checker_entries_barrier_2_io_y_hw = dcache_pma_checker_entries_barrier_2_io_y_hw;
    assign dcache__pma_checker_entries_barrier_2_io_y_hx = dcache_pma_checker_entries_barrier_2_io_y_hx;
    assign dcache__pma_checker_entries_barrier_2_io_y_hr = dcache_pma_checker_entries_barrier_2_io_y_hr;
    assign dcache__pma_checker_entries_barrier_2_io_y_pw = dcache_pma_checker_entries_barrier_2_io_y_pw;
    assign dcache__pma_checker_entries_barrier_2_io_y_px = dcache_pma_checker_entries_barrier_2_io_y_px;
    assign dcache__pma_checker_entries_barrier_2_io_y_pr = dcache_pma_checker_entries_barrier_2_io_y_pr;
    assign dcache__pma_checker_entries_barrier_2_io_y_ppp = dcache_pma_checker_entries_barrier_2_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_2_io_y_pal = dcache_pma_checker_entries_barrier_2_io_y_pal;
    assign dcache__pma_checker_entries_barrier_2_io_y_paa = dcache_pma_checker_entries_barrier_2_io_y_paa;
    assign dcache__pma_checker_entries_barrier_2_io_y_eff = dcache_pma_checker_entries_barrier_2_io_y_eff;
    assign dcache__pma_checker_entries_barrier_2_io_y_c = dcache_pma_checker_entries_barrier_2_io_y_c;
    assign dcache_pma_checker_entries_barrier_3_io_x_u = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_ae_ptw = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_ae_final = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_ae_stage2 = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_pf = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_gf = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_sw = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_sx = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_sr = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_hw = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_hx = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_hr = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_pw = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_px = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_pr = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_ppp = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_pal = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_paa = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_eff = 1'h0;
    assign dcache_pma_checker_entries_barrier_3_io_x_c = 1'h0;
    assign dcache__pma_checker_entries_barrier_3_io_y_u = dcache_pma_checker_entries_barrier_3_io_y_u;
    assign dcache__pma_checker_entries_barrier_3_io_y_ae_ptw = dcache_pma_checker_entries_barrier_3_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_3_io_y_ae_final = dcache_pma_checker_entries_barrier_3_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_3_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_3_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_3_io_y_pf = dcache_pma_checker_entries_barrier_3_io_y_pf;
    assign dcache__pma_checker_entries_barrier_3_io_y_gf = dcache_pma_checker_entries_barrier_3_io_y_gf;
    assign dcache__pma_checker_entries_barrier_3_io_y_sw = dcache_pma_checker_entries_barrier_3_io_y_sw;
    assign dcache__pma_checker_entries_barrier_3_io_y_sx = dcache_pma_checker_entries_barrier_3_io_y_sx;
    assign dcache__pma_checker_entries_barrier_3_io_y_sr = dcache_pma_checker_entries_barrier_3_io_y_sr;
    assign dcache__pma_checker_entries_barrier_3_io_y_hw = dcache_pma_checker_entries_barrier_3_io_y_hw;
    assign dcache__pma_checker_entries_barrier_3_io_y_hx = dcache_pma_checker_entries_barrier_3_io_y_hx;
    assign dcache__pma_checker_entries_barrier_3_io_y_hr = dcache_pma_checker_entries_barrier_3_io_y_hr;
    assign dcache__pma_checker_entries_barrier_3_io_y_pw = dcache_pma_checker_entries_barrier_3_io_y_pw;
    assign dcache__pma_checker_entries_barrier_3_io_y_px = dcache_pma_checker_entries_barrier_3_io_y_px;
    assign dcache__pma_checker_entries_barrier_3_io_y_pr = dcache_pma_checker_entries_barrier_3_io_y_pr;
    assign dcache__pma_checker_entries_barrier_3_io_y_ppp = dcache_pma_checker_entries_barrier_3_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_3_io_y_pal = dcache_pma_checker_entries_barrier_3_io_y_pal;
    assign dcache__pma_checker_entries_barrier_3_io_y_paa = dcache_pma_checker_entries_barrier_3_io_y_paa;
    assign dcache__pma_checker_entries_barrier_3_io_y_eff = dcache_pma_checker_entries_barrier_3_io_y_eff;
    assign dcache__pma_checker_entries_barrier_3_io_y_c = dcache_pma_checker_entries_barrier_3_io_y_c;
    assign dcache_pma_checker_entries_barrier_4_io_x_u = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_ae_ptw = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_ae_final = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_ae_stage2 = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_pf = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_gf = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_sw = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_sx = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_sr = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_hw = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_hx = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_hr = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_pw = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_px = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_pr = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_ppp = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_pal = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_paa = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_eff = 1'h0;
    assign dcache_pma_checker_entries_barrier_4_io_x_c = 1'h0;
    assign dcache__pma_checker_entries_barrier_4_io_y_u = dcache_pma_checker_entries_barrier_4_io_y_u;
    assign dcache__pma_checker_entries_barrier_4_io_y_ae_ptw = dcache_pma_checker_entries_barrier_4_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_4_io_y_ae_final = dcache_pma_checker_entries_barrier_4_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_4_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_4_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_4_io_y_pf = dcache_pma_checker_entries_barrier_4_io_y_pf;
    assign dcache__pma_checker_entries_barrier_4_io_y_gf = dcache_pma_checker_entries_barrier_4_io_y_gf;
    assign dcache__pma_checker_entries_barrier_4_io_y_sw = dcache_pma_checker_entries_barrier_4_io_y_sw;
    assign dcache__pma_checker_entries_barrier_4_io_y_sx = dcache_pma_checker_entries_barrier_4_io_y_sx;
    assign dcache__pma_checker_entries_barrier_4_io_y_sr = dcache_pma_checker_entries_barrier_4_io_y_sr;
    assign dcache__pma_checker_entries_barrier_4_io_y_hw = dcache_pma_checker_entries_barrier_4_io_y_hw;
    assign dcache__pma_checker_entries_barrier_4_io_y_hx = dcache_pma_checker_entries_barrier_4_io_y_hx;
    assign dcache__pma_checker_entries_barrier_4_io_y_hr = dcache_pma_checker_entries_barrier_4_io_y_hr;
    assign dcache__pma_checker_entries_barrier_4_io_y_pw = dcache_pma_checker_entries_barrier_4_io_y_pw;
    assign dcache__pma_checker_entries_barrier_4_io_y_px = dcache_pma_checker_entries_barrier_4_io_y_px;
    assign dcache__pma_checker_entries_barrier_4_io_y_pr = dcache_pma_checker_entries_barrier_4_io_y_pr;
    assign dcache__pma_checker_entries_barrier_4_io_y_ppp = dcache_pma_checker_entries_barrier_4_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_4_io_y_pal = dcache_pma_checker_entries_barrier_4_io_y_pal;
    assign dcache__pma_checker_entries_barrier_4_io_y_paa = dcache_pma_checker_entries_barrier_4_io_y_paa;
    assign dcache__pma_checker_entries_barrier_4_io_y_eff = dcache_pma_checker_entries_barrier_4_io_y_eff;
    assign dcache__pma_checker_entries_barrier_4_io_y_c = dcache_pma_checker_entries_barrier_4_io_y_c;
    assign dcache_pma_checker_entries_barrier_5_io_x_u = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_ae_ptw = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_ae_final = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_ae_stage2 = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_pf = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_gf = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_sw = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_sx = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_sr = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_hw = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_hx = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_hr = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_pw = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_px = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_pr = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_ppp = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_pal = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_paa = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_eff = 1'h0;
    assign dcache_pma_checker_entries_barrier_5_io_x_c = 1'h0;
    assign dcache__pma_checker_entries_barrier_5_io_y_u = dcache_pma_checker_entries_barrier_5_io_y_u;
    assign dcache__pma_checker_entries_barrier_5_io_y_ae_ptw = dcache_pma_checker_entries_barrier_5_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_5_io_y_ae_final = dcache_pma_checker_entries_barrier_5_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_5_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_5_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_5_io_y_pf = dcache_pma_checker_entries_barrier_5_io_y_pf;
    assign dcache__pma_checker_entries_barrier_5_io_y_gf = dcache_pma_checker_entries_barrier_5_io_y_gf;
    assign dcache__pma_checker_entries_barrier_5_io_y_sw = dcache_pma_checker_entries_barrier_5_io_y_sw;
    assign dcache__pma_checker_entries_barrier_5_io_y_sx = dcache_pma_checker_entries_barrier_5_io_y_sx;
    assign dcache__pma_checker_entries_barrier_5_io_y_sr = dcache_pma_checker_entries_barrier_5_io_y_sr;
    assign dcache__pma_checker_entries_barrier_5_io_y_hw = dcache_pma_checker_entries_barrier_5_io_y_hw;
    assign dcache__pma_checker_entries_barrier_5_io_y_hx = dcache_pma_checker_entries_barrier_5_io_y_hx;
    assign dcache__pma_checker_entries_barrier_5_io_y_hr = dcache_pma_checker_entries_barrier_5_io_y_hr;
      
    wire dcache_lfsr_prng_clock;
    wire dcache_lfsr_prng_reset;
    wire dcache_lfsr_prng_io_increment;
    wire dcache_lfsr_prng_io_out_0;
    wire dcache_lfsr_prng_io_out_1;
    wire dcache_lfsr_prng_io_out_2;
    wire dcache_lfsr_prng_io_out_3;
    wire dcache_lfsr_prng_io_out_4;
    wire dcache_lfsr_prng_io_out_5;
    wire dcache_lfsr_prng_io_out_6;
    wire dcache_lfsr_prng_io_out_7;
    wire dcache_lfsr_prng_io_out_8;
    wire dcache_lfsr_prng_io_out_9;
    wire dcache_lfsr_prng_io_out_10;
    wire dcache_lfsr_prng_io_out_11;
    wire dcache_lfsr_prng_io_out_12;
    wire dcache_lfsr_prng_io_out_13;
    wire dcache_lfsr_prng_io_out_14;
    wire dcache_lfsr_prng_io_out_15;

    reg dcache_lfsr_prng_state_0 ; 
    reg dcache_lfsr_prng_state_1 ; 
    reg dcache_lfsr_prng_state_2 ; 
    reg dcache_lfsr_prng_state_3 ; 
    reg dcache_lfsr_prng_state_4 ; 
    reg dcache_lfsr_prng_state_5 ; 
    reg dcache_lfsr_prng_state_6 ; 
    reg dcache_lfsr_prng_state_7 ; 
    reg dcache_lfsr_prng_state_8 ; 
    reg dcache_lfsr_prng_state_9 ; 
    reg dcache_lfsr_prng_state_10 ; 
    reg dcache_lfsr_prng_state_11 ; 
    reg dcache_lfsr_prng_state_12 ; 
    reg dcache_lfsr_prng_state_13 ; 
    reg dcache_lfsr_prng_state_14 ; 
    reg dcache_lfsr_prng_state_15 ; 
  always @( posedge  dcache_lfsr_prng_clock )
         begin 
             if ( dcache_lfsr_prng_reset )
                 begin  
                     dcache_lfsr_prng_state_0  <=1'h1; 
                     dcache_lfsr_prng_state_1  <=1'h0; 
                     dcache_lfsr_prng_state_2  <=1'h0; 
                     dcache_lfsr_prng_state_3  <=1'h0; 
                     dcache_lfsr_prng_state_4  <=1'h0; 
                     dcache_lfsr_prng_state_5  <=1'h0; 
                     dcache_lfsr_prng_state_6  <=1'h0; 
                     dcache_lfsr_prng_state_7  <=1'h0; 
                     dcache_lfsr_prng_state_8  <=1'h0; 
                     dcache_lfsr_prng_state_9  <=1'h0; 
                     dcache_lfsr_prng_state_10  <=1'h0; 
                     dcache_lfsr_prng_state_11  <=1'h0; 
                     dcache_lfsr_prng_state_12  <=1'h0; 
                     dcache_lfsr_prng_state_13  <=1'h0; 
                     dcache_lfsr_prng_state_14  <=1'h0; 
                     dcache_lfsr_prng_state_15  <=1'h0;
                 end 
              else 
                 if ( dcache_lfsr_prng_io_increment )
                     begin  
                         dcache_lfsr_prng_state_0  <= dcache_lfsr_prng_state_15 ^ dcache_lfsr_prng_state_13 ^ dcache_lfsr_prng_state_12 ^ dcache_lfsr_prng_state_10 ; 
                         dcache_lfsr_prng_state_1  <= dcache_lfsr_prng_state_0 ; 
                         dcache_lfsr_prng_state_2  <= dcache_lfsr_prng_state_1 ; 
                         dcache_lfsr_prng_state_3  <= dcache_lfsr_prng_state_2 ; 
                         dcache_lfsr_prng_state_4  <= dcache_lfsr_prng_state_3 ; 
                         dcache_lfsr_prng_state_5  <= dcache_lfsr_prng_state_4 ; 
                         dcache_lfsr_prng_state_6  <= dcache_lfsr_prng_state_5 ; 
                         dcache_lfsr_prng_state_7  <= dcache_lfsr_prng_state_6 ; 
                         dcache_lfsr_prng_state_8  <= dcache_lfsr_prng_state_7 ; 
                         dcache_lfsr_prng_state_9  <= dcache_lfsr_prng_state_8 ; 
                         dcache_lfsr_prng_state_10  <= dcache_lfsr_prng_state_9 ; 
                         dcache_lfsr_prng_state_11  <= dcache_lfsr_prng_state_10 ; 
                         dcache_lfsr_prng_state_12  <= dcache_lfsr_prng_state_11 ; 
                         dcache_lfsr_prng_state_13  <= dcache_lfsr_prng_state_12 ; 
                         dcache_lfsr_prng_state_14  <= dcache_lfsr_prng_state_13 ; 
                         dcache_lfsr_prng_state_15  <= dcache_lfsr_prng_state_14 ;
                     end 
         end
  assign  dcache_lfsr_prng_io_out_0 = dcache_lfsr_prng_state_0 ; 
  assign  dcache_lfsr_prng_io_out_1 = dcache_lfsr_prng_state_1 ; 
  assign  dcache_lfsr_prng_io_out_2 = dcache_lfsr_prng_state_2 ; 
  assign  dcache_lfsr_prng_io_out_3 = dcache_lfsr_prng_state_3 ; 
  assign  dcache_lfsr_prng_io_out_4 = dcache_lfsr_prng_state_4 ; 
  assign  dcache_lfsr_prng_io_out_5 = dcache_lfsr_prng_state_5 ; 
  assign  dcache_lfsr_prng_io_out_6 = dcache_lfsr_prng_state_6 ; 
  assign  dcache_lfsr_prng_io_out_7 = dcache_lfsr_prng_state_7 ; 
  assign  dcache_lfsr_prng_io_out_8 = dcache_lfsr_prng_state_8 ; 
  assign  dcache_lfsr_prng_io_out_9 = dcache_lfsr_prng_state_9 ; 
  assign  dcache_lfsr_prng_io_out_10 = dcache_lfsr_prng_state_10 ; 
  assign  dcache_lfsr_prng_io_out_11 = dcache_lfsr_prng_state_11 ; 
  assign  dcache_lfsr_prng_io_out_12 = dcache_lfsr_prng_state_12 ; 
  assign  dcache_lfsr_prng_io_out_13 = dcache_lfsr_prng_state_13 ; 
  assign  dcache_lfsr_prng_io_out_14 = dcache_lfsr_prng_state_14 ; 
  assign  dcache_lfsr_prng_io_out_15 = dcache_lfsr_prng_state_15 ;
    assign dcache_lfsr_prng_clock = dcache_clock;
    assign dcache_lfsr_prng_reset = dcache_reset;
    assign dcache_lfsr_prng_io_increment = dcache_replace;
    assign dcache__lfsr_prng_io_out_0 = dcache_lfsr_prng_io_out_0;
    assign dcache__lfsr_prng_io_out_1 = dcache_lfsr_prng_io_out_1;
    assign dcache__lfsr_prng_io_out_2 = dcache_lfsr_prng_io_out_2;
    assign dcache__lfsr_prng_io_out_3 = dcache_lfsr_prng_io_out_3;
    assign dcache__lfsr_prng_io_out_4 = dcache_lfsr_prng_io_out_4;
    assign dcache__lfsr_prng_io_out_5 = dcache_lfsr_prng_io_out_5;
    assign dcache__lfsr_prng_io_out_6 = dcache_lfsr_prng_io_out_6;
    assign dcache__lfsr_prng_io_out_7 = dcache_lfsr_prng_io_out_7;
    assign dcache__lfsr_prng_io_out_8 = dcache_lfsr_prng_io_out_8;
    assign dcache__lfsr_prng_io_out_9 = dcache_lfsr_prng_io_out_9;
    assign dcache__lfsr_prng_io_out_10 = dcache_lfsr_prng_io_out_10;
    assign dcache__lfsr_prng_io_out_11 = dcache_lfsr_prng_io_out_11;
    assign dcache__lfsr_prng_io_out_12 = dcache_lfsr_prng_io_out_12;
    assign dcache__lfsr_prng_io_out_13 = dcache_lfsr_prng_io_out_13;
    assign dcache__lfsr_prng_io_out_14 = dcache_lfsr_prng_io_out_14;
    assign dcache__lfsr_prng_io_out_15 = dcache_lfsr_prng_io_out_15;
      
    wire dcache_data_clock;
    wire dcache_data_io_req_valid;
    wire[13:0] dcache_data_io_req_bits_addr;
    wire dcache_data_io_req_bits_write;
    wire[31:0] dcache_data_io_req_bits_wdata;
    wire[3:0] dcache_data_io_req_bits_eccMask;
    wire[31:0] dcache_data_io_resp_0;

    wire dcache_data_data_arrays_0_rdata_data_en ; 
    wire dcache_data_data_arrays_0_rdata_MPORT_en ; 
    wire[31:0] dcache_data__data_arrays_0_ext_RW0_rdata ; 
    wire[31:0] dcache_data_wWords_0 = dcache_data_io_req_bits_wdata ; 
    wire dcache_data_rdata_valid = dcache_data_io_req_valid ; 
    wire dcache_data_eccMask_0 = dcache_data_io_req_bits_eccMask [0]; 
    wire dcache_data_eccMask_1 = dcache_data_io_req_bits_eccMask [1]; 
    wire dcache_data_eccMask_2 = dcache_data_io_req_bits_eccMask [2]; 
    wire dcache_data_eccMask_3 = dcache_data_io_req_bits_eccMask [3]; 
    wire[11:0] dcache_data_addr = dcache_data_io_req_bits_addr [13:2]; 
    wire[7:0] dcache_data_rdata_wData_0 ; 
    wire[7:0] dcache_data_rdata_wData_1 ; 
    wire[7:0] dcache_data_rdata_wData_2 ; 
    wire[7:0] dcache_data_rdata_wData_3 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_en = dcache_data_rdata_valid & dcache_data_io_req_bits_write ; 
  assign  dcache_data_rdata_wData_0 = dcache_data_wWords_0 [7:0]; 
  assign  dcache_data_rdata_wData_1 = dcache_data_wWords_0 [15:8]; 
  assign  dcache_data_rdata_wData_2 = dcache_data_wWords_0 [23:16]; 
  assign  dcache_data_rdata_wData_3 = dcache_data_wWords_0 [31:24]; 
  assign  dcache_data_data_arrays_0_rdata_data_en = dcache_data_rdata_valid &~ dcache_data_io_req_bits_write ; 
    wire[15:0] dcache_data_rdata_lo = dcache_data__data_arrays_0_ext_RW0_rdata [15:0]; 
    wire[15:0] dcache_data_rdata_hi = dcache_data__data_arrays_0_ext_RW0_rdata [31:16]; 
    wire[31:0] dcache_data_rdata_0_0 ={ dcache_data_rdata_hi , dcache_data_rdata_lo };  
    wire[11:0] dcache_data_data_arrays_0_ext_RW0_addr;
    wire dcache_data_data_arrays_0_ext_RW0_en;
    wire dcache_data_data_arrays_0_ext_RW0_clk;
    wire dcache_data_data_arrays_0_ext_RW0_wmode;
    wire[31:0] dcache_data_data_arrays_0_ext_RW0_wdata;
    wire[31:0] dcache_data_data_arrays_0_ext_RW0_rdata;
    wire[3:0] dcache_data_data_arrays_0_ext_RW0_wmask;

    reg[31:0] dcache_data_data_arrays_0_ext_Memory [0:4095]; reg[11:0] dcache_data_data_arrays_0_ext__RW0_raddr_d0 ; 
    reg dcache_data_data_arrays_0_ext__RW0_ren_d0 ; 
    reg dcache_data_data_arrays_0_ext__RW0_rmode_d0 ; 
  always @( posedge  dcache_data_data_arrays_0_ext_RW0_clk )
         begin  
             dcache_data_data_arrays_0_ext__RW0_raddr_d0  <= dcache_data_data_arrays_0_ext_RW0_addr ; 
             dcache_data_data_arrays_0_ext__RW0_ren_d0  <= dcache_data_data_arrays_0_ext_RW0_en ; 
             dcache_data_data_arrays_0_ext__RW0_rmode_d0  <= dcache_data_data_arrays_0_ext_RW0_wmode ;
             if ( dcache_data_data_arrays_0_ext_RW0_en & dcache_data_data_arrays_0_ext_RW0_wmask [0]& dcache_data_data_arrays_0_ext_RW0_wmode ) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_RW0_addr ][32'h0+:8]<= dcache_data_data_arrays_0_ext_RW0_wdata [7:0];
             if ( dcache_data_data_arrays_0_ext_RW0_en & dcache_data_data_arrays_0_ext_RW0_wmask [1]& dcache_data_data_arrays_0_ext_RW0_wmode ) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_RW0_addr ][32'h8+:8]<= dcache_data_data_arrays_0_ext_RW0_wdata [15:8];
             if ( dcache_data_data_arrays_0_ext_RW0_en & dcache_data_data_arrays_0_ext_RW0_wmask [2]& dcache_data_data_arrays_0_ext_RW0_wmode ) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_RW0_addr ][32'h10+:8]<= dcache_data_data_arrays_0_ext_RW0_wdata [23:16];
             if ( dcache_data_data_arrays_0_ext_RW0_en & dcache_data_data_arrays_0_ext_RW0_wmask [3]& dcache_data_data_arrays_0_ext_RW0_wmode ) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_RW0_addr ][32'h18+:8]<= dcache_data_data_arrays_0_ext_RW0_wdata [31:24];
         end
  assign  dcache_data_data_arrays_0_ext_RW0_rdata = dcache_data_data_arrays_0_ext__RW0_ren_d0 &~ dcache_data_data_arrays_0_ext__RW0_rmode_d0  ?  dcache_data_data_arrays_0_ext_Memory [ dcache_data_data_arrays_0_ext__RW0_raddr_d0 ]:32'bx;
    assign dcache_data_data_arrays_0_ext_RW0_addr = dcache_data_addr;
    assign dcache_data_data_arrays_0_ext_RW0_en = dcache_data_data_arrays_0_rdata_data_en|dcache_data_data_arrays_0_rdata_MPORT_en;
    assign dcache_data_data_arrays_0_ext_RW0_clk = dcache_data_clock;
    assign dcache_data_data_arrays_0_ext_RW0_wmode = dcache_data_io_req_bits_write;
    assign dcache_data_data_arrays_0_ext_RW0_wdata = {dcache_data_rdata_wData_3,dcache_data_rdata_wData_2,dcache_data_rdata_wData_1,dcache_data_rdata_wData_0};
    assign dcache_data__data_arrays_0_ext_RW0_rdata = dcache_data_data_arrays_0_ext_RW0_rdata;
    assign dcache_data_data_arrays_0_ext_RW0_wmask = {dcache_data_eccMask_3,dcache_data_eccMask_2,dcache_data_eccMask_1,dcache_data_eccMask_0};
     
  assign  dcache_data_io_resp_0 = dcache_data_rdata_0_0 ;
    assign dcache_data_clock = dcache_clock;
    assign dcache_data_io_req_valid = dcache_dataArb_io_out_valid;
    assign dcache_data_io_req_bits_addr = dcache__GEN_46 ? dcache__dataArb_io_in_0_bits_wordMask_wordMask_T:dcache_dataArb_io_in_3_bits_addr;
    assign dcache_data_io_req_bits_write = (dcache_dataArb_io_in_0_valid|dcache_dataArb_io_in_1_valid&dcache__GEN)&dcache_pstore_drain;
    assign dcache_data_io_req_bits_wdata = {dcache_dataArb_io_in_0_bits_wdata_hi,dcache_dataArb_io_in_0_bits_wdata_lo};
    assign dcache_data_io_req_bits_eccMask = dcache__GEN_46 ? dcache_dataArb_io_in_1_bits_eccMask:4'hF;
    assign dcache_s1_all_data_ways_0 = dcache_data_io_resp_0;
      
    wire[3:0] dcache_amoalus_0_io_mask;
    wire[4:0] dcache_amoalus_0_io_cmd;
    wire[31:0] dcache_amoalus_0_io_lhs;
    wire[31:0] dcache_amoalus_0_io_rhs;
    wire[31:0] dcache_amoalus_0_io_out_unmasked;

    wire[31:0] dcache_amoalus_0_adder_out_mask =32'hFFFFFFFF; 
    wire[3:0] dcache_amoalus_0_less_signed_mask =4'h2; 
    wire dcache_amoalus_0_max = dcache_amoalus_0_io_cmd ==5'hD| dcache_amoalus_0_io_cmd ==5'hF; 
    wire dcache_amoalus_0_min = dcache_amoalus_0_io_cmd ==5'hC| dcache_amoalus_0_io_cmd ==5'hE; 
    wire dcache_amoalus_0_add = dcache_amoalus_0_io_cmd ==5'h8; 
    wire dcache_amoalus_0__logic_xor_T_1 = dcache_amoalus_0_io_cmd ==5'hA; 
    wire dcache_amoalus_0_logic_and = dcache_amoalus_0__logic_xor_T_1 | dcache_amoalus_0_io_cmd ==5'hB; 
    wire dcache_amoalus_0_logic_xor = dcache_amoalus_0_io_cmd ==5'h9| dcache_amoalus_0__logic_xor_T_1 ; 
    wire[31:0] dcache_amoalus_0_adder_out = dcache_amoalus_0_io_lhs + dcache_amoalus_0_io_rhs ; 
    wire dcache_amoalus_0_less_signed =~( dcache_amoalus_0_io_cmd [1]); 
    wire dcache_amoalus_0_less = dcache_amoalus_0_io_lhs [31]== dcache_amoalus_0_io_rhs [31] ?  dcache_amoalus_0_io_lhs < dcache_amoalus_0_io_rhs : dcache_amoalus_0_less_signed  ?  dcache_amoalus_0_io_lhs [31]: dcache_amoalus_0_io_rhs [31]; 
    wire[31:0] dcache_amoalus_0_minmax =( dcache_amoalus_0_less  ?  dcache_amoalus_0_min : dcache_amoalus_0_max ) ?  dcache_amoalus_0_io_lhs : dcache_amoalus_0_io_rhs ; 
    wire[31:0] dcache_amoalus_0_logic_0 =( dcache_amoalus_0_logic_and  ?  dcache_amoalus_0_io_lhs & dcache_amoalus_0_io_rhs :32'h0)|( dcache_amoalus_0_logic_xor  ?  dcache_amoalus_0_io_lhs ^ dcache_amoalus_0_io_rhs :32'h0); 
    wire[31:0] dcache_amoalus_0_out = dcache_amoalus_0_add  ?  dcache_amoalus_0_adder_out : dcache_amoalus_0_logic_and | dcache_amoalus_0_logic_xor  ?  dcache_amoalus_0_logic_0 : dcache_amoalus_0_minmax ; 
    wire[15:0] dcache_amoalus_0_wmask_lo ={{8{ dcache_amoalus_0_io_mask [1]}},{8{ dcache_amoalus_0_io_mask [0]}}}; 
    wire[15:0] dcache_amoalus_0_wmask_hi ={{8{ dcache_amoalus_0_io_mask [3]}},{8{ dcache_amoalus_0_io_mask [2]}}}; 
    wire[31:0] dcache_amoalus_0_wmask ={ dcache_amoalus_0_wmask_hi , dcache_amoalus_0_wmask_lo }; 
  assign  dcache_amoalus_0_io_out_unmasked = dcache_amoalus_0_out ;
    assign dcache_amoalus_0_io_mask = dcache_pstore1_mask;
    assign dcache_amoalus_0_io_cmd = dcache_pstore1_cmd;
    assign dcache_amoalus_0_io_lhs = dcache_s2_data_word;
    assign dcache_amoalus_0_io_rhs = dcache_pstore1_data;
    assign dcache__amoalus_0_io_out_unmasked = dcache_amoalus_0_io_out_unmasked;
     
  assign  dcache_auto_out_a_valid = dcache_nodeOut_a_valid ; 
  assign  dcache_auto_out_a_bits_opcode = dcache_nodeOut_a_bits_opcode ; 
  assign  dcache_auto_out_a_bits_param = dcache_nodeOut_a_bits_param ; 
  assign  dcache_auto_out_a_bits_size = dcache_nodeOut_a_bits_size ; 
  assign  dcache_auto_out_a_bits_address = dcache_nodeOut_a_bits_address ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_bufferable = dcache_nodeOut_a_bits_user_amba_prot_bufferable ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_modifiable = dcache_nodeOut_a_bits_user_amba_prot_modifiable ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_readalloc = dcache_nodeOut_a_bits_user_amba_prot_readalloc ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_writealloc = dcache_nodeOut_a_bits_user_amba_prot_writealloc ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_privileged = dcache_nodeOut_a_bits_user_amba_prot_privileged ; 
  assign  dcache_auto_out_a_bits_mask = dcache_nodeOut_a_bits_mask ; 
  assign  dcache_auto_out_a_bits_data = dcache_nodeOut_a_bits_data ; 
  assign  dcache_auto_out_d_ready = dcache_nodeOut_d_ready ; 
  assign  dcache_io_cpu_req_ready = dcache__io_cpu_req_ready_output ; 
  assign  dcache_io_cpu_s2_nack = dcache__io_cpu_s2_nack_output ; 
  assign  dcache_io_cpu_resp_valid = dcache_s2_valid_hit_pre_data_ecc | dcache_doUncachedResp ; 
  assign  dcache_io_cpu_resp_bits_addr = dcache_doUncachedResp  ?  dcache_s2_uncached_resp_addr : dcache_s2_req_addr ; 
  assign  dcache_io_cpu_resp_bits_tag = dcache_s2_req_tag ; 
  assign  dcache_io_cpu_resp_bits_cmd = dcache_s2_req_cmd ; 
  assign  dcache_io_cpu_resp_bits_size = dcache_s2_req_size ; 
  assign  dcache_io_cpu_resp_bits_signed = dcache_s2_req_signed ; 
  assign  dcache_io_cpu_resp_bits_dprv = dcache_s2_req_dprv ; 
  assign  dcache_io_cpu_resp_bits_dv = dcache_s2_req_dv ; 
  assign  dcache_io_cpu_resp_bits_data ={ dcache_size ==2'h0 ? {24{ dcache_s2_req_signed & dcache_io_cpu_resp_bits_data_zeroed_1 [7]}}:{ dcache_size ==2'h1 ? {16{ dcache_s2_req_signed & dcache_io_cpu_resp_bits_data_zeroed [15]}}: dcache_s2_data_word_possibly_uncached [31:16], dcache_io_cpu_resp_bits_data_zeroed [15:8]}, dcache_io_cpu_resp_bits_data_zeroed_1 }; 
  assign  dcache_io_cpu_resp_bits_mask = dcache_s2_req_mask ; 
  assign  dcache_io_cpu_resp_bits_replay = dcache_doUncachedResp ; 
  assign  dcache_io_cpu_resp_bits_has_data = dcache_s2_read ; 
  assign  dcache_io_cpu_resp_bits_data_word_bypass = dcache_s2_data_word_possibly_uncached ; 
  assign  dcache_io_cpu_resp_bits_data_raw = dcache_s2_data_word ; 
  assign  dcache_io_cpu_resp_bits_store_data = dcache_pstore1_data ; 
  assign  dcache_io_cpu_replay_next = dcache__io_cpu_replay_next_output ; 
  assign  dcache_io_cpu_s2_xcpt_ma_ld = dcache__io_cpu_s2_xcpt_ma_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_ma_st = dcache__io_cpu_s2_xcpt_ma_st_output ; 
  assign  dcache_io_cpu_s2_xcpt_pf_ld = dcache__io_cpu_s2_xcpt_pf_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_pf_st = dcache__io_cpu_s2_xcpt_pf_st_output ; 
  assign  dcache_io_cpu_s2_xcpt_ae_ld = dcache__io_cpu_s2_xcpt_ae_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_ae_st = dcache__io_cpu_s2_xcpt_ae_st_output ; 
  assign  dcache_io_cpu_ordered =~( dcache_s1_valid &~ dcache_s1_req_no_xcpt | dcache_s2_valid &~ dcache_s2_req_no_xcpt | dcache_cached_grant_wait | dcache_uncachedInFlight_0 ); 
  assign  dcache_io_cpu_perf_grant = dcache_nodeOut_d_valid & dcache_d_last ; 
  assign  dcache_io_ptw_req_bits_bits_addr =20'h0; 
  assign  dcache_io_ptw_req_bits_bits_need_gpa =1'h0; 
  assign  dcache_io_ptw_req_bits_bits_vstage1 =1'h0; 
  assign  dcache_io_ptw_req_bits_bits_stage2 =1'h0;
    assign dcache_clock = clock;
    assign dcache_reset = reset;
    assign dcache_auto_hart_id_sink_in = broadcast_x1_nodeOut;
    assign dcache_auto_out_a_ready = widget_nodeIn_a_ready;
    assign widget_nodeIn_a_valid = dcache_auto_out_a_valid;
    assign widget_nodeIn_a_bits_opcode = dcache_auto_out_a_bits_opcode;
    assign widget_nodeIn_a_bits_param = dcache_auto_out_a_bits_param;
    assign widget_nodeIn_a_bits_size = dcache_auto_out_a_bits_size;
    assign widget_nodeIn_a_bits_address = dcache_auto_out_a_bits_address;
    assign widget_nodeIn_a_bits_user_amba_prot_bufferable = dcache_auto_out_a_bits_user_amba_prot_bufferable;
    assign widget_nodeIn_a_bits_user_amba_prot_modifiable = dcache_auto_out_a_bits_user_amba_prot_modifiable;
    assign widget_nodeIn_a_bits_user_amba_prot_readalloc = dcache_auto_out_a_bits_user_amba_prot_readalloc;
    assign widget_nodeIn_a_bits_user_amba_prot_writealloc = dcache_auto_out_a_bits_user_amba_prot_writealloc;
    assign widget_nodeIn_a_bits_user_amba_prot_privileged = dcache_auto_out_a_bits_user_amba_prot_privileged;
    assign widget_nodeIn_a_bits_mask = dcache_auto_out_a_bits_mask;
    assign widget_nodeIn_a_bits_data = dcache_auto_out_a_bits_data;
    assign widget_nodeIn_d_ready = dcache_auto_out_d_ready;
    assign dcache_auto_out_d_valid = widget_nodeIn_d_valid;
    assign dcache_auto_out_d_bits_opcode = widget_nodeIn_d_bits_opcode;
    assign dcache_auto_out_d_bits_param = widget_nodeIn_d_bits_param;
    assign dcache_auto_out_d_bits_size = widget_nodeIn_d_bits_size;
    assign dcache_auto_out_d_bits_sink = widget_nodeIn_d_bits_sink;
    assign dcache_auto_out_d_bits_denied = widget_nodeIn_d_bits_denied;
    assign dcache_auto_out_d_bits_data = widget_nodeIn_d_bits_data;
    assign dcache_auto_out_d_bits_corrupt = widget_nodeIn_d_bits_corrupt;
    assign _dcache_io_cpu_req_ready = dcache_io_cpu_req_ready;
    assign dcache_io_cpu_req_valid = _dcacheArb_io_mem_req_valid;
    assign dcache_io_cpu_req_bits_addr = _dcacheArb_io_mem_req_bits_addr;
    assign dcache_io_cpu_req_bits_tag = _dcacheArb_io_mem_req_bits_tag;
    assign dcache_io_cpu_req_bits_cmd = _dcacheArb_io_mem_req_bits_cmd;
    assign dcache_io_cpu_req_bits_size = _dcacheArb_io_mem_req_bits_size;
    assign dcache_io_cpu_req_bits_signed = _dcacheArb_io_mem_req_bits_signed;
    assign dcache_io_cpu_req_bits_dprv = _dcacheArb_io_mem_req_bits_dprv;
    assign dcache_io_cpu_req_bits_dv = _dcacheArb_io_mem_req_bits_dv;
    assign dcache_io_cpu_req_bits_phys = _dcacheArb_io_mem_req_bits_phys;
    assign dcache_io_cpu_req_bits_no_xcpt = _dcacheArb_io_mem_req_bits_no_xcpt;
    assign dcache_io_cpu_s1_kill = _dcacheArb_io_mem_s1_kill;
    assign dcache_io_cpu_s1_data_data = _dcacheArb_io_mem_s1_data_data;
    assign dcache_io_cpu_s1_data_mask = _dcacheArb_io_mem_s1_data_mask;
    assign _dcache_io_cpu_s2_nack = dcache_io_cpu_s2_nack;
    assign _dcache_io_cpu_resp_valid = dcache_io_cpu_resp_valid;
    assign _dcache_io_cpu_resp_bits_tag = dcache_io_cpu_resp_bits_tag;
    assign _dcache_io_cpu_resp_bits_data = dcache_io_cpu_resp_bits_data;
    assign _dcache_io_cpu_resp_bits_replay = dcache_io_cpu_resp_bits_replay;
    assign _dcache_io_cpu_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data;
    assign _dcache_io_cpu_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass;
    assign _dcache_io_cpu_resp_bits_data_raw = dcache_io_cpu_resp_bits_data_raw;
    assign _dcache_io_cpu_replay_next = dcache_io_cpu_replay_next;
    assign _dcache_io_cpu_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld;
    assign _dcache_io_cpu_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st;
    assign _dcache_io_cpu_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld;
    assign _dcache_io_cpu_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st;
    assign _dcache_io_cpu_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld;
    assign _dcache_io_cpu_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st;
    assign _dcache_io_cpu_ordered = dcache_io_cpu_ordered;
    assign _dcache_io_cpu_perf_grant = dcache_io_cpu_perf_grant;
    assign _dcache_io_ptw_req_bits_bits_addr = dcache_io_ptw_req_bits_bits_addr;
    assign _dcache_io_ptw_req_bits_bits_need_gpa = dcache_io_ptw_req_bits_bits_need_gpa;
    assign _dcache_io_ptw_req_bits_bits_vstage1 = dcache_io_ptw_req_bits_bits_vstage1;
    assign _dcache_io_ptw_req_bits_bits_stage2 = dcache_io_ptw_req_bits_bits_stage2;
    assign dcache_io_ptw_resp_bits_ae_ptw = _ptw_io_requestor_0_resp_bits_ae_ptw;
    assign dcache_io_ptw_resp_bits_ae_final = _ptw_io_requestor_0_resp_bits_ae_final;
    assign dcache_io_ptw_resp_bits_pf = _ptw_io_requestor_0_resp_bits_pf;
    assign dcache_io_ptw_resp_bits_gf = _ptw_io_requestor_0_resp_bits_gf;
    assign dcache_io_ptw_resp_bits_hr = _ptw_io_requestor_0_resp_bits_hr;
    assign dcache_io_ptw_resp_bits_hw = _ptw_io_requestor_0_resp_bits_hw;
    assign dcache_io_ptw_resp_bits_hx = _ptw_io_requestor_0_resp_bits_hx;
    assign dcache_io_ptw_resp_bits_pte_ppn = _ptw_io_requestor_0_resp_bits_pte_ppn;
    assign dcache_io_ptw_resp_bits_pte_d = _ptw_io_requestor_0_resp_bits_pte_d;
    assign dcache_io_ptw_resp_bits_pte_a = _ptw_io_requestor_0_resp_bits_pte_a;
    assign dcache_io_ptw_resp_bits_pte_g = _ptw_io_requestor_0_resp_bits_pte_g;
    assign dcache_io_ptw_resp_bits_pte_u = _ptw_io_requestor_0_resp_bits_pte_u;
    assign dcache_io_ptw_resp_bits_pte_x = _ptw_io_requestor_0_resp_bits_pte_x;
    assign dcache_io_ptw_resp_bits_pte_w = _ptw_io_requestor_0_resp_bits_pte_w;
    assign dcache_io_ptw_resp_bits_pte_r = _ptw_io_requestor_0_resp_bits_pte_r;
    assign dcache_io_ptw_resp_bits_pte_v = _ptw_io_requestor_0_resp_bits_pte_v;
    assign dcache_io_ptw_resp_bits_gpa_is_pte = _ptw_io_requestor_0_resp_bits_gpa_is_pte;
    assign dcache_io_ptw_status_debug = _ptw_io_requestor_0_status_debug;
    assign dcache_io_ptw_pmp_0_cfg_l = _ptw_io_requestor_0_pmp_0_cfg_l;
    assign dcache_io_ptw_pmp_0_cfg_a = _ptw_io_requestor_0_pmp_0_cfg_a;
    assign dcache_io_ptw_pmp_0_cfg_x = _ptw_io_requestor_0_pmp_0_cfg_x;
    assign dcache_io_ptw_pmp_0_cfg_w = _ptw_io_requestor_0_pmp_0_cfg_w;
    assign dcache_io_ptw_pmp_0_cfg_r = _ptw_io_requestor_0_pmp_0_cfg_r;
    assign dcache_io_ptw_pmp_0_addr = _ptw_io_requestor_0_pmp_0_addr;
    assign dcache_io_ptw_pmp_0_mask = _ptw_io_requestor_0_pmp_0_mask;
    assign dcache_io_ptw_pmp_1_cfg_l = _ptw_io_requestor_0_pmp_1_cfg_l;
    assign dcache_io_ptw_pmp_1_cfg_a = _ptw_io_requestor_0_pmp_1_cfg_a;
    assign dcache_io_ptw_pmp_1_cfg_x = _ptw_io_requestor_0_pmp_1_cfg_x;
    assign dcache_io_ptw_pmp_1_cfg_w = _ptw_io_requestor_0_pmp_1_cfg_w;
    assign dcache_io_ptw_pmp_1_cfg_r = _ptw_io_requestor_0_pmp_1_cfg_r;
    assign dcache_io_ptw_pmp_1_addr = _ptw_io_requestor_0_pmp_1_addr;
    assign dcache_io_ptw_pmp_1_mask = _ptw_io_requestor_0_pmp_1_mask;
    assign dcache_io_ptw_pmp_2_cfg_l = _ptw_io_requestor_0_pmp_2_cfg_l;
    assign dcache_io_ptw_pmp_2_cfg_a = _ptw_io_requestor_0_pmp_2_cfg_a;
    assign dcache_io_ptw_pmp_2_cfg_x = _ptw_io_requestor_0_pmp_2_cfg_x;
    assign dcache_io_ptw_pmp_2_cfg_w = _ptw_io_requestor_0_pmp_2_cfg_w;
    assign dcache_io_ptw_pmp_2_cfg_r = _ptw_io_requestor_0_pmp_2_cfg_r;
    assign dcache_io_ptw_pmp_2_addr = _ptw_io_requestor_0_pmp_2_addr;
    assign dcache_io_ptw_pmp_2_mask = _ptw_io_requestor_0_pmp_2_mask;
    assign dcache_io_ptw_pmp_3_cfg_l = _ptw_io_requestor_0_pmp_3_cfg_l;
    assign dcache_io_ptw_pmp_3_cfg_a = _ptw_io_requestor_0_pmp_3_cfg_a;
    assign dcache_io_ptw_pmp_3_cfg_x = _ptw_io_requestor_0_pmp_3_cfg_x;
    assign dcache_io_ptw_pmp_3_cfg_w = _ptw_io_requestor_0_pmp_3_cfg_w;
    assign dcache_io_ptw_pmp_3_cfg_r = _ptw_io_requestor_0_pmp_3_cfg_r;
    assign dcache_io_ptw_pmp_3_addr = _ptw_io_requestor_0_pmp_3_addr;
    assign dcache_io_ptw_pmp_3_mask = _ptw_io_requestor_0_pmp_3_mask;
    assign dcache_io_ptw_pmp_4_cfg_l = _ptw_io_requestor_0_pmp_4_cfg_l;
    assign dcache_io_ptw_pmp_4_cfg_a = _ptw_io_requestor_0_pmp_4_cfg_a;
    assign dcache_io_ptw_pmp_4_cfg_x = _ptw_io_requestor_0_pmp_4_cfg_x;
    assign dcache_io_ptw_pmp_4_cfg_w = _ptw_io_requestor_0_pmp_4_cfg_w;
    assign dcache_io_ptw_pmp_4_cfg_r = _ptw_io_requestor_0_pmp_4_cfg_r;
    assign dcache_io_ptw_pmp_4_addr = _ptw_io_requestor_0_pmp_4_addr;
    assign dcache_io_ptw_pmp_4_mask = _ptw_io_requestor_0_pmp_4_mask;
    assign dcache_io_ptw_pmp_5_cfg_l = _ptw_io_requestor_0_pmp_5_cfg_l;
    assign dcache_io_ptw_pmp_5_cfg_a = _ptw_io_requestor_0_pmp_5_cfg_a;
    assign dcache_io_ptw_pmp_5_cfg_x = _ptw_io_requestor_0_pmp_5_cfg_x;
    assign dcache_io_ptw_pmp_5_cfg_w = _ptw_io_requestor_0_pmp_5_cfg_w;
    assign dcache_io_ptw_pmp_5_cfg_r = _ptw_io_requestor_0_pmp_5_cfg_r;
    assign dcache_io_ptw_pmp_5_addr = _ptw_io_requestor_0_pmp_5_addr;
    assign dcache_io_ptw_pmp_5_mask = _ptw_io_requestor_0_pmp_5_mask;
    assign dcache_io_ptw_pmp_6_cfg_l = _ptw_io_requestor_0_pmp_6_cfg_l;
    assign dcache_io_ptw_pmp_6_cfg_a = _ptw_io_requestor_0_pmp_6_cfg_a;
    assign dcache_io_ptw_pmp_6_cfg_x = _ptw_io_requestor_0_pmp_6_cfg_x;
    assign dcache_io_ptw_pmp_6_cfg_w = _ptw_io_requestor_0_pmp_6_cfg_w;
    assign dcache_io_ptw_pmp_6_cfg_r = _ptw_io_requestor_0_pmp_6_cfg_r;
    assign dcache_io_ptw_pmp_6_addr = _ptw_io_requestor_0_pmp_6_addr;
    assign dcache_io_ptw_pmp_6_mask = _ptw_io_requestor_0_pmp_6_mask;
    assign dcache_io_ptw_pmp_7_cfg_l = _ptw_io_requestor_0_pmp_7_cfg_l;
    assign dcache_io_ptw_pmp_7_cfg_a = _ptw_io_requestor_0_pmp_7_cfg_a;
    assign dcache_io_ptw_pmp_7_cfg_x = _ptw_io_requestor_0_pmp_7_cfg_x;
    assign dcache_io_ptw_pmp_7_cfg_w = _ptw_io_requestor_0_pmp_7_cfg_w;
    assign dcache_io_ptw_pmp_7_cfg_r = _ptw_io_requestor_0_pmp_7_cfg_r;
    assign dcache_io_ptw_pmp_7_addr = _ptw_io_requestor_0_pmp_7_addr;
    assign dcache_io_ptw_pmp_7_mask = _ptw_io_requestor_0_pmp_7_mask;
    
  wire frontend_clock;
    wire frontend_reset;
    wire frontend_auto_icache_master_out_a_ready;
    wire frontend_auto_icache_master_out_a_valid;
    wire[31:0] frontend_auto_icache_master_out_a_bits_address;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_readalloc;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_writealloc;
    wire frontend_auto_icache_master_out_d_valid;
    wire[2:0] frontend_auto_icache_master_out_d_bits_opcode;
    wire[1:0] frontend_auto_icache_master_out_d_bits_param;
    wire[3:0] frontend_auto_icache_master_out_d_bits_size;
    wire frontend_auto_icache_master_out_d_bits_sink;
    wire frontend_auto_icache_master_out_d_bits_denied;
    wire[31:0] frontend_auto_icache_master_out_d_bits_data;
    wire frontend_auto_icache_master_out_d_bits_corrupt;
    wire frontend_io_cpu_might_request;
    wire frontend_io_cpu_req_valid;
    wire[31:0] frontend_io_cpu_req_bits_pc;
    wire frontend_io_cpu_req_bits_speculative;
    wire frontend_io_cpu_sfence_valid;
    wire frontend_io_cpu_resp_ready;
    wire frontend_io_cpu_resp_valid;
    wire[1:0] frontend_io_cpu_resp_bits_btb_cfiType;
    wire frontend_io_cpu_resp_bits_btb_taken;
    wire[1:0] frontend_io_cpu_resp_bits_btb_mask;
    wire frontend_io_cpu_resp_bits_btb_bridx;
    wire[31:0] frontend_io_cpu_resp_bits_btb_target;
    wire frontend_io_cpu_resp_bits_btb_entry;
    wire[7:0] frontend_io_cpu_resp_bits_btb_bht_history;
    wire frontend_io_cpu_resp_bits_btb_bht_value;
    wire[31:0] frontend_io_cpu_resp_bits_pc;
    wire[31:0] frontend_io_cpu_resp_bits_data;
    wire[1:0] frontend_io_cpu_resp_bits_mask;
    wire frontend_io_cpu_resp_bits_xcpt_pf_inst;
    wire frontend_io_cpu_resp_bits_xcpt_gf_inst;
    wire frontend_io_cpu_resp_bits_xcpt_ae_inst;
    wire frontend_io_cpu_resp_bits_replay;
    wire frontend_io_cpu_gpa_valid;
    wire[31:0] frontend_io_cpu_gpa_bits;
    wire frontend_io_cpu_btb_update_valid;
    wire frontend_io_cpu_bht_update_valid;
    wire frontend_io_cpu_flush_icache;
    wire frontend_io_cpu_progress;
    wire frontend_io_ptw_req_bits_valid;
    wire[19:0] frontend_io_ptw_req_bits_bits_addr;
    wire frontend_io_ptw_req_bits_bits_need_gpa;
    wire frontend_io_ptw_req_bits_bits_vstage1;
    wire frontend_io_ptw_req_bits_bits_stage2;
    wire frontend_io_ptw_resp_bits_ae_ptw;
    wire frontend_io_ptw_resp_bits_ae_final;
    wire frontend_io_ptw_resp_bits_pf;
    wire frontend_io_ptw_resp_bits_gf;
    wire frontend_io_ptw_resp_bits_hr;
    wire frontend_io_ptw_resp_bits_hw;
    wire frontend_io_ptw_resp_bits_hx;
    wire[43:0] frontend_io_ptw_resp_bits_pte_ppn;
    wire frontend_io_ptw_resp_bits_pte_d;
    wire frontend_io_ptw_resp_bits_pte_a;
    wire frontend_io_ptw_resp_bits_pte_g;
    wire frontend_io_ptw_resp_bits_pte_u;
    wire frontend_io_ptw_resp_bits_pte_x;
    wire frontend_io_ptw_resp_bits_pte_w;
    wire frontend_io_ptw_resp_bits_pte_r;
    wire frontend_io_ptw_resp_bits_pte_v;
    wire frontend_io_ptw_resp_bits_gpa_is_pte;
    wire frontend_io_ptw_status_debug;
    wire frontend_io_ptw_pmp_0_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_0_cfg_a;
    wire frontend_io_ptw_pmp_0_cfg_x;
    wire frontend_io_ptw_pmp_0_cfg_w;
    wire frontend_io_ptw_pmp_0_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_0_addr;
    wire[31:0] frontend_io_ptw_pmp_0_mask;
    wire frontend_io_ptw_pmp_1_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_1_cfg_a;
    wire frontend_io_ptw_pmp_1_cfg_x;
    wire frontend_io_ptw_pmp_1_cfg_w;
    wire frontend_io_ptw_pmp_1_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_1_addr;
    wire[31:0] frontend_io_ptw_pmp_1_mask;
    wire frontend_io_ptw_pmp_2_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_2_cfg_a;
    wire frontend_io_ptw_pmp_2_cfg_x;
    wire frontend_io_ptw_pmp_2_cfg_w;
    wire frontend_io_ptw_pmp_2_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_2_addr;
    wire[31:0] frontend_io_ptw_pmp_2_mask;
    wire frontend_io_ptw_pmp_3_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_3_cfg_a;
    wire frontend_io_ptw_pmp_3_cfg_x;
    wire frontend_io_ptw_pmp_3_cfg_w;
    wire frontend_io_ptw_pmp_3_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_3_addr;
    wire[31:0] frontend_io_ptw_pmp_3_mask;
    wire frontend_io_ptw_pmp_4_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_4_cfg_a;
    wire frontend_io_ptw_pmp_4_cfg_x;
    wire frontend_io_ptw_pmp_4_cfg_w;
    wire frontend_io_ptw_pmp_4_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_4_addr;
    wire[31:0] frontend_io_ptw_pmp_4_mask;
    wire frontend_io_ptw_pmp_5_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_5_cfg_a;
    wire frontend_io_ptw_pmp_5_cfg_x;
    wire frontend_io_ptw_pmp_5_cfg_w;
    wire frontend_io_ptw_pmp_5_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_5_addr;
    wire[31:0] frontend_io_ptw_pmp_5_mask;
    wire frontend_io_ptw_pmp_6_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_6_cfg_a;
    wire frontend_io_ptw_pmp_6_cfg_x;
    wire frontend_io_ptw_pmp_6_cfg_w;
    wire frontend_io_ptw_pmp_6_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_6_addr;
    wire[31:0] frontend_io_ptw_pmp_6_mask;
    wire frontend_io_ptw_pmp_7_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_7_cfg_a;
    wire frontend_io_ptw_pmp_7_cfg_x;
    wire frontend_io_ptw_pmp_7_cfg_w;
    wire frontend_io_ptw_pmp_7_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_7_addr;
    wire[31:0] frontend_io_ptw_pmp_7_mask;
    wire[31:0] frontend_io_ptw_customCSRs_csrs_0_value;

    wire frontend__fq_io_enq_valid_T_6 ; 
    wire[31:0] frontend__tlb_io_resp_paddr ; 
    wire[31:0] frontend__tlb_io_resp_gpa ; 
    wire frontend__tlb_io_resp_pf_ld ; 
    wire frontend__tlb_io_resp_pf_inst ; 
    wire frontend__tlb_io_resp_ae_ld ; 
    wire frontend__tlb_io_resp_ae_inst ; 
    wire frontend__tlb_io_resp_ma_ld ; 
    wire frontend__tlb_io_resp_cacheable ; 
    wire frontend__tlb_io_resp_prefetchable ; 
    wire frontend__fq_io_enq_ready ; 
    wire[4:0] frontend__fq_io_mask ; 
    wire frontend__icache_io_resp_valid ; 
    wire[31:0] frontend__icache_io_resp_bits_data ; 
    wire frontend__icache_io_resp_bits_ae ; 
    wire frontend_s2_redirect = frontend_io_cpu_req_valid ; 
    wire frontend_s2_btb_taken =1'h0; 
    wire frontend_predicted_taken =1'h0; 
    wire frontend_clock_en =1'h1; 
    wire[31:0] frontend_resetVectorSinkNodeIn =32'h10040; 
    reg frontend_s1_valid ; 
    reg frontend_s2_valid ; 
    wire frontend_s0_fq_has_space =~( frontend__fq_io_mask [2])|~( frontend__fq_io_mask [3])&(~ frontend_s1_valid |~ frontend_s2_valid )|~( frontend__fq_io_mask [4])&~ frontend_s1_valid &~ frontend_s2_valid ; 
    wire frontend_s0_valid = frontend_io_cpu_req_valid | frontend_s0_fq_has_space ; reg[31:0] frontend_s1_pc ; 
    reg frontend_s1_speculative ; reg[31:0] frontend_s2_pc ; reg[31:0] frontend_s2_tlb_resp_paddr ; reg[31:0] frontend_s2_tlb_resp_gpa ; 
    reg frontend_s2_tlb_resp_pf_ld ; 
    reg frontend_s2_tlb_resp_pf_inst ; 
    reg frontend_s2_tlb_resp_ae_ld ; 
    reg frontend_s2_tlb_resp_ae_inst ; 
    reg frontend_s2_tlb_resp_ma_ld ; 
    reg frontend_s2_tlb_resp_cacheable ; 
    reg frontend_s2_tlb_resp_prefetchable ; 
    wire frontend_s2_xcpt = frontend_s2_tlb_resp_ae_inst | frontend_s2_tlb_resp_pf_inst ; 
    reg frontend_s2_speculative ; 
    wire[31:0] frontend_s1_base_pc ={ frontend_s1_pc [31:2],2'h0}; 
    wire[31:0] frontend_ntpc = frontend_s1_base_pc +32'h4; 
    wire[31:0] frontend_predicted_npc = frontend_ntpc ; 
    reg frontend_s2_replay_REG ; 
    wire frontend_s2_replay = frontend_s2_valid &~( frontend__fq_io_enq_ready & frontend__fq_io_enq_valid_T_6 )| frontend_s2_replay_REG ; 
    wire[31:0] frontend_npc = frontend_s2_replay  ?  frontend_s2_pc : frontend_predicted_npc ; 
    wire frontend_s0_speculative = frontend_s1_speculative | frontend_s2_valid &~ frontend_s2_speculative ; reg[1:0] frontend_recent_progress_counter ; 
    wire frontend_recent_progress =| frontend_recent_progress_counter ; 
    wire frontend_s2_kill_speculative_tlb_refill = frontend_s2_speculative &~ frontend_recent_progress ; 
    wire frontend_s2_can_speculatively_refill = frontend_s2_tlb_resp_cacheable &~( frontend_io_ptw_customCSRs_csrs_0_value [3]); 
    wire frontend__icache_io_s2_kill_T_2 = frontend_s2_speculative &~ frontend_s2_can_speculatively_refill | frontend_s2_xcpt ; 
    reg frontend_fq_io_enq_valid_REG ; 
  assign  frontend__fq_io_enq_valid_T_6 = frontend_fq_io_enq_valid_REG & frontend_s2_valid &( frontend__icache_io_resp_valid | frontend__icache_io_s2_kill_T_2 ); 
    wire[31:0] frontend__io_cpu_npc_T_3 ={ frontend_io_cpu_req_valid  ?  frontend_io_cpu_req_bits_pc [31:1]: frontend_npc [31:1],1'h0}; 
    wire[2:0] frontend__fq_io_enq_bits_mask_T_1 =3'h3<< frontend_s2_pc [1]; 
  always @( posedge  frontend_clock )
         begin 
             if (~ frontend_reset &~(~( frontend_io_cpu_req_valid | frontend_io_cpu_sfence_valid | frontend_io_cpu_flush_icache | frontend_io_cpu_bht_update_valid | frontend_io_cpu_btb_update_valid )| frontend_io_cpu_might_request ))
                 begin 
                     if (1)$error("Assertion failed\n    at Frontend.scala:92 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n");
                     if (1)$fatal;
                 end 
             if (~ frontend_reset & frontend_s2_speculative & frontend_io_ptw_customCSRs_csrs_0_value [3]&~ frontend__icache_io_s2_kill_T_2 )
                 begin 
                     if (1)$error("Assertion failed\n    at Frontend.scala:190 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n");
                     if (1)$fatal;
                 end 
         end
    reg frontend_gpa_valid ; reg[31:0] frontend_gpa ; 
  always @( posedge  frontend_clock )
         begin  
             frontend_s1_valid  <= frontend_s0_valid ; 
             frontend_s1_pc  <= frontend__io_cpu_npc_T_3 ;
             if ( frontend_io_cpu_req_valid ) 
                 frontend_s1_speculative  <= frontend_io_cpu_req_bits_speculative ;
              else 
                 if ( frontend_s2_replay ) 
                     frontend_s1_speculative  <= frontend_s2_speculative ;
                  else  
                     frontend_s1_speculative  <= frontend_s0_speculative ;
             if ( frontend_s2_replay )
                 begin 
                 end 
              else 
                 begin  
                     frontend_s2_tlb_resp_paddr  <= frontend__tlb_io_resp_paddr ; 
                     frontend_s2_tlb_resp_gpa  <= frontend__tlb_io_resp_gpa ; 
                     frontend_s2_tlb_resp_pf_ld  <= frontend__tlb_io_resp_pf_ld ; 
                     frontend_s2_tlb_resp_pf_inst  <= frontend__tlb_io_resp_pf_inst ; 
                     frontend_s2_tlb_resp_ae_ld  <= frontend__tlb_io_resp_ae_ld ; 
                     frontend_s2_tlb_resp_ae_inst  <= frontend__tlb_io_resp_ae_inst ; 
                     frontend_s2_tlb_resp_ma_ld  <= frontend__tlb_io_resp_ma_ld ; 
                     frontend_s2_tlb_resp_cacheable  <= frontend__tlb_io_resp_cacheable ; 
                     frontend_s2_tlb_resp_prefetchable  <= frontend__tlb_io_resp_prefetchable ;
                 end  
             frontend_fq_io_enq_valid_REG  <= frontend_s1_valid ;
             if ( frontend_reset )
                 begin  
                     frontend_s2_valid  <=1'h0; 
                     frontend_s2_pc  <=32'h10040; 
                     frontend_s2_speculative  <=1'h0; 
                     frontend_s2_replay_REG  <=1'h1; 
                     frontend_recent_progress_counter  <=2'h3;
                 end 
              else 
                 begin  
                     frontend_s2_valid  <=~ frontend_s2_replay &~ frontend_s2_redirect ;
                     if ( frontend_s2_replay )
                         begin 
                         end 
                      else 
                         begin  
                             frontend_s2_pc  <= frontend_s1_pc ; 
                             frontend_s2_speculative  <= frontend_s1_speculative ;
                         end  
                     frontend_s2_replay_REG  <= frontend_s2_replay &~ frontend_s0_valid ;
                     if ( frontend_io_cpu_progress ) 
                         frontend_recent_progress_counter  <=2'h3;
                 end 
             if ( frontend_io_cpu_req_valid ) 
                 frontend_gpa_valid  <=1'h0;
         end
    wire frontend_icache_clock;
    wire frontend_icache_reset;
    wire frontend_icache_auto_master_out_a_ready;
    wire frontend_icache_auto_master_out_a_valid;
    wire[31:0] frontend_icache_auto_master_out_a_bits_address;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_readalloc;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_writealloc;
    wire frontend_icache_auto_master_out_d_valid;
    wire[2:0] frontend_icache_auto_master_out_d_bits_opcode;
    wire[1:0] frontend_icache_auto_master_out_d_bits_param;
    wire[3:0] frontend_icache_auto_master_out_d_bits_size;
    wire frontend_icache_auto_master_out_d_bits_sink;
    wire frontend_icache_auto_master_out_d_bits_denied;
    wire[31:0] frontend_icache_auto_master_out_d_bits_data;
    wire frontend_icache_auto_master_out_d_bits_corrupt;
    wire frontend_icache_io_req_valid;
    wire[31:0] frontend_icache_io_req_bits_addr;
    wire[31:0] frontend_icache_io_s1_paddr;
    wire[31:0] frontend_icache_io_s2_vaddr;
    wire frontend_icache_io_s1_kill;
    wire frontend_icache_io_s2_kill;
    wire frontend_icache_io_s2_cacheable;
    wire frontend_icache_io_resp_valid;
    wire[31:0] frontend_icache_io_resp_bits_data;
    wire frontend_icache_io_resp_bits_ae;
    wire frontend_icache_io_invalidate;

    wire frontend_icache_readEnable ; 
    wire frontend_icache_readEnable_0 ; 
    wire[5:0] frontend_icache__tag_rdata_T_4 ; 
    wire frontend_icache__io_req_ready_T_2 ; 
    wire[20:0] frontend_icache__tag_array_0_ext_RW0_rdata ; 
    wire frontend_icache_masterNodeOut_a_ready = frontend_icache_auto_master_out_a_ready ; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_readalloc = frontend_icache_io_s2_cacheable ; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_writealloc = frontend_icache_io_s2_cacheable ; 
    wire frontend_icache_masterNodeOut_d_valid = frontend_icache_auto_master_out_d_valid ; 
    wire[2:0] frontend_icache_masterNodeOut_d_bits_opcode = frontend_icache_auto_master_out_d_bits_opcode ; 
    wire[1:0] frontend_icache_masterNodeOut_d_bits_param = frontend_icache_auto_master_out_d_bits_param ; 
    wire[3:0] frontend_icache_masterNodeOut_d_bits_size = frontend_icache_auto_master_out_d_bits_size ; 
    wire frontend_icache_masterNodeOut_d_bits_sink = frontend_icache_auto_master_out_d_bits_sink ; 
    wire frontend_icache_masterNodeOut_d_bits_denied = frontend_icache_auto_master_out_d_bits_denied ; 
    wire[31:0] frontend_icache_masterNodeOut_d_bits_data = frontend_icache_auto_master_out_d_bits_data ; 
    wire frontend_icache_masterNodeOut_d_bits_corrupt = frontend_icache_auto_master_out_d_bits_corrupt ; 
    wire frontend_icache_invalidate = frontend_icache_io_invalidate ; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_bufferable =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_modifiable =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_privileged =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_secure =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_fetch =1'h1; 
    wire frontend_icache_masterNodeOut_d_ready =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_1 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_size_1 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_2 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_3 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_4 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_5 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_source =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_corrupt =1'h0; 
    wire frontend_icache_masterNodeOut_d_bits_source =1'h0; 
    wire frontend_icache_s1_tag_disparity_0 =1'h0; 
    wire frontend_icache_scratchpadHit =1'h0; 
    wire frontend_icache_way =1'h0; 
    wire frontend_icache_s1s2_full_word_write =1'h0; 
    wire frontend_icache_s1_dont_read =1'h0; 
    wire frontend_icache_s2_tag_disparity =1'h0; 
    wire frontend_icache_s2_disparity =1'h0; 
    wire frontend_icache_s1_scratchpad_hit =1'h0; 
    wire frontend_icache_s2_report_uncorrectable_error =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_source =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_bufferable =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_modifiable =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_readalloc =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_writealloc =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_privileged =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_secure =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_fetch =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_corrupt =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH_shiftAmount =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_size =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_bit =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 =1'h0; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_param =3'h0; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_a_param =3'h0; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_opcode =3'h4; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_a_opcode =3'h4; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_size =4'h6; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_a_size =4'h6; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_mask =4'hF; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_a_mask =4'hF; 
    wire[31:0] frontend_icache_masterNodeOut_a_bits_data =32'h0; 
    wire[31:0] frontend_icache_masterNodeOut_a_bits_a_data =32'h0; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_lo =2'h3; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_hi =2'h3; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH =2'h1; 
    wire frontend_icache_s2_request_refill ; 
    wire[31:0] frontend_icache_masterNodeOut_a_bits_a_address ; 
    wire[31:0] frontend_icache_data = frontend_icache_masterNodeOut_d_bits_data ; 
    wire frontend_icache_s0_valid = frontend_icache__io_req_ready_T_2 & frontend_icache_io_req_valid ; 
    wire frontend_icache_s0_ren = frontend_icache_s0_valid ; 
    reg frontend_icache_s1_valid ; 
    wire frontend_icache_s1_clk_en = frontend_icache_s1_valid ; reg[31:0] frontend_icache_s1_vaddr ; 
    wire frontend_icache_tagMatch ; 
    wire frontend_icache_s1_tag_hit_0 ; 
    wire frontend_icache_s1_hit = frontend_icache_s1_tag_hit_0 ; 
    reg frontend_icache_s2_valid ; 
    reg frontend_icache_s2_hit ; 
    reg frontend_icache_invalidated ; 
    reg frontend_icache_refill_valid ; 
    wire frontend_icache_masterNodeOut_a_valid ; 
    wire frontend_icache_refill_fire = frontend_icache_masterNodeOut_a_ready & frontend_icache_masterNodeOut_a_valid ; 
    wire frontend_icache_s2_miss = frontend_icache_s2_valid &~ frontend_icache_s2_hit &~ frontend_icache_io_s2_kill ; 
    wire frontend_icache_s1_can_request_refill =~( frontend_icache_s2_miss | frontend_icache_refill_valid ); 
    reg frontend_icache_s2_request_refill_REG ; 
  assign  frontend_icache_s2_request_refill = frontend_icache_s2_miss & frontend_icache_s2_request_refill_REG ; 
  assign  frontend_icache_masterNodeOut_a_valid = frontend_icache_s2_request_refill ; reg[31:0] frontend_icache_refill_paddr ; reg[31:0] frontend_icache_refill_vaddr ; 
    wire[19:0] frontend_icache_refill_tag = frontend_icache_refill_paddr [31:12]; 
    wire[5:0] frontend_icache_refill_idx = frontend_icache_refill_paddr [11:6]; 
    wire frontend_icache_refill_one_beat_opdata = frontend_icache_masterNodeOut_d_bits_opcode [0]; 
    wire frontend_icache_beats1_opdata = frontend_icache_masterNodeOut_d_bits_opcode [0]; 
    wire frontend_icache_refill_one_beat = frontend_icache_masterNodeOut_d_valid & frontend_icache_refill_one_beat_opdata ; 
  assign  frontend_icache__io_req_ready_T_2 =~ frontend_icache_refill_one_beat ; 
    wire[26:0] frontend_icache__beats1_decode_T_1 =27'hFFF<< frontend_icache_masterNodeOut_d_bits_size ; 
    wire[9:0] frontend_icache_beats1_decode =~( frontend_icache__beats1_decode_T_1 [11:2]); 
    wire[9:0] frontend_icache_beats1 = frontend_icache_beats1_opdata  ?  frontend_icache_beats1_decode :10'h0; reg[9:0] frontend_icache_counter ; 
    wire[9:0] frontend_icache_counter1 = frontend_icache_counter -10'h1; 
    wire frontend_icache_first = frontend_icache_counter ==10'h0; 
    wire frontend_icache_last = frontend_icache_counter ==10'h1| frontend_icache_beats1 ==10'h0; 
    wire frontend_icache_d_done = frontend_icache_last & frontend_icache_masterNodeOut_d_valid ; 
    wire[9:0] frontend_icache_refill_cnt = frontend_icache_beats1 &~ frontend_icache_counter1 ; 
    wire frontend_icache_refill_done = frontend_icache_refill_one_beat & frontend_icache_d_done ; 
  assign  frontend_icache__tag_rdata_T_4 = frontend_icache_io_req_bits_addr [11:6]; 
  assign  frontend_icache_readEnable_0 =~ frontend_icache_refill_done & frontend_icache_s0_valid ; 
    reg frontend_icache_accruedRefillError ; 
    wire frontend_icache_refillError = frontend_icache_masterNodeOut_d_bits_corrupt |(| frontend_icache_refill_cnt )& frontend_icache_accruedRefillError ; 
    wire[20:0] frontend_icache_enc_tag ={ frontend_icache_refillError , frontend_icache_refill_tag }; reg[63:0] frontend_icache_vb_array ; 
    wire[5:0] frontend_icache_s1_idx = frontend_icache_io_s1_paddr [11:6]; 
    wire[19:0] frontend_icache_s1_tag = frontend_icache_io_s1_paddr [31:12]; 
    wire[63:0] frontend_icache__s1_vb_T_1 = frontend_icache_vb_array >> frontend_icache_s1_idx ; 
    wire frontend_icache_s1_vb = frontend_icache__s1_vb_T_1 [0]; 
    wire frontend_icache_tl_error = frontend_icache__tag_array_0_ext_RW0_rdata [20]; 
    wire[19:0] frontend_icache_tag = frontend_icache__tag_array_0_ext_RW0_rdata [19:0]; 
  assign  frontend_icache_tagMatch = frontend_icache_s1_vb & frontend_icache_tag == frontend_icache_s1_tag ; 
  assign  frontend_icache_s1_tag_hit_0 = frontend_icache_tagMatch ; 
    wire frontend_icache_s1_tl_error_0 = frontend_icache_tagMatch & frontend_icache_tl_error ; 
    wire frontend_icache_wen ; 
  assign  frontend_icache_wen = frontend_icache_refill_one_beat &~ frontend_icache_invalidated ; 
    wire[9:0] frontend_icache_mem_idx = frontend_icache_refill_one_beat  ? { frontend_icache_refill_idx ,4'h0}| frontend_icache_refill_cnt : frontend_icache_io_req_bits_addr [11:2]; 
  assign  frontend_icache_readEnable =~ frontend_icache_wen & frontend_icache_s0_ren ; 
    reg frontend_icache_s2_tag_hit_0 ; 
    wire[10:0] frontend_icache_s2_scratchpad_word_addr_hi ={1'h0, frontend_icache_io_s2_vaddr [11:2]}; 
    wire[12:0] frontend_icache_s2_scratchpad_word_addr ={ frontend_icache_s2_scratchpad_word_addr_hi ,2'h0}; reg[31:0] frontend_icache_s2_dout_0 ; 
    reg frontend_icache_s2_tl_error ; 
  assign  frontend_icache_masterNodeOut_a_bits_a_address ={ frontend_icache_refill_paddr [31:6],6'h0}; 
    wire frontend_icache_masterNodeOut_a_bits_legal ={ frontend_icache_refill_paddr [31:30], frontend_icache_refill_paddr [27], frontend_icache_refill_paddr [25], frontend_icache_refill_paddr [16],~( frontend_icache_refill_paddr [13])}==6'h0|{ frontend_icache_refill_paddr [31:30], frontend_icache_refill_paddr [27], frontend_icache_refill_paddr [25], frontend_icache_refill_paddr [16], frontend_icache_refill_paddr [13]}==6'h0|{ frontend_icache_refill_paddr [31:30], frontend_icache_refill_paddr [27], frontend_icache_refill_paddr [25],~( frontend_icache_refill_paddr [16])}==5'h0|{ frontend_icache_refill_paddr [31:30], frontend_icache_refill_paddr [27],~( frontend_icache_refill_paddr [25]), frontend_icache_refill_paddr [16]}==5'h0|{ frontend_icache_refill_paddr [31:30],~( frontend_icache_refill_paddr [27])}==3'h0|{ frontend_icache_refill_paddr [31],~( frontend_icache_refill_paddr [30])}==2'h0|{ frontend_icache_refill_paddr [31:30]^2'h2, frontend_icache_refill_paddr [27], frontend_icache_refill_paddr [25], frontend_icache_refill_paddr [16]}==5'h0; 
    wire[31:0] frontend_icache_masterNodeOut_a_bits_address = frontend_icache_masterNodeOut_a_bits_a_address ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_1 = frontend_icache_masterNodeOut_a_bits_a_mask_bit ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_nbit =~ frontend_icache_masterNodeOut_a_bits_a_mask_bit ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq = frontend_icache_masterNodeOut_a_bits_a_mask_nbit ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_nbit_1 =~ frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_2 = frontend_icache_masterNodeOut_a_bits_a_mask_eq & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_3 = frontend_icache_masterNodeOut_a_bits_a_mask_eq & frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_4 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_1 & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_5 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_1 & frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 ; 
    wire[127:0] frontend_icache__vb_array_T_3 =128'h1<< frontend_icache_refill_idx ; 
    wire[31:0] frontend_icache_s1_dout_0 ; 
  always @( posedge  frontend_icache_clock )
         begin 
             if ( frontend_icache_reset )
                 begin  
                     frontend_icache_s1_valid  <=1'h0; 
                     frontend_icache_s2_valid  <=1'h0; 
                     frontend_icache_refill_valid  <=1'h0; 
                     frontend_icache_counter  <=10'h0; 
                     frontend_icache_vb_array  <=64'h0;
                 end 
              else 
                 begin  
                     frontend_icache_s1_valid  <= frontend_icache_s0_valid ; 
                     frontend_icache_s2_valid  <= frontend_icache_s1_valid &~ frontend_icache_io_s1_kill ; 
                     frontend_icache_refill_valid  <=~ frontend_icache_refill_done &( frontend_icache_refill_fire | frontend_icache_refill_valid );
                     if ( frontend_icache_masterNodeOut_d_valid )
                         begin 
                             if ( frontend_icache_first ) 
                                 frontend_icache_counter  <= frontend_icache_beats1 ;
                              else  
                                 frontend_icache_counter  <= frontend_icache_counter1 ;
                         end 
                     if ( frontend_icache_invalidate ) 
                         frontend_icache_vb_array  <=64'h0;
                      else 
                         if ( frontend_icache_refill_one_beat ) 
                             frontend_icache_vb_array  <= frontend_icache_refill_done &~ frontend_icache_invalidated  ?  frontend_icache_vb_array | frontend_icache__vb_array_T_3 [63:0]:~(~ frontend_icache_vb_array | frontend_icache__vb_array_T_3 [63:0]);
                 end 
             if ( frontend_icache_s0_valid ) 
                 frontend_icache_s1_vaddr  <= frontend_icache_io_req_bits_addr ; 
             frontend_icache_s2_hit  <= frontend_icache_s1_hit ; 
             frontend_icache_invalidated  <= frontend_icache_refill_valid &( frontend_icache_invalidate | frontend_icache_invalidated ); 
             frontend_icache_s2_request_refill_REG  <= frontend_icache_s1_can_request_refill ;
             if ( frontend_icache_s1_valid & frontend_icache_s1_can_request_refill )
                 begin  
                     frontend_icache_refill_paddr  <= frontend_icache_io_s1_paddr ; 
                     frontend_icache_refill_vaddr  <= frontend_icache_s1_vaddr ;
                 end 
             if ( frontend_icache_refill_one_beat ) 
                 frontend_icache_accruedRefillError  <= frontend_icache_refillError ;
             if ( frontend_icache_s1_clk_en )
                 begin  
                     frontend_icache_s2_tag_hit_0  <= frontend_icache_s1_tag_hit_0 ; 
                     frontend_icache_s2_dout_0  <= frontend_icache_s1_dout_0 ; 
                     frontend_icache_s2_tl_error  <= frontend_icache_s1_tl_error_0 ;
                 end 
         end
    wire[5:0] frontend_icache_tag_array_0_ext_RW0_addr;
    wire frontend_icache_tag_array_0_ext_RW0_en;
    wire frontend_icache_tag_array_0_ext_RW0_clk;
    wire frontend_icache_tag_array_0_ext_RW0_wmode;
    wire[20:0] frontend_icache_tag_array_0_ext_RW0_wdata;
    wire[20:0] frontend_icache_tag_array_0_ext_RW0_rdata;

    reg[20:0] frontend_icache_tag_array_0_ext_Memory [0:63]; reg[5:0] frontend_icache_tag_array_0_ext__RW0_raddr_d0 ; 
    reg frontend_icache_tag_array_0_ext__RW0_ren_d0 ; 
    reg frontend_icache_tag_array_0_ext__RW0_rmode_d0 ; 
  always @( posedge  frontend_icache_tag_array_0_ext_RW0_clk )
         begin  
             frontend_icache_tag_array_0_ext__RW0_raddr_d0  <= frontend_icache_tag_array_0_ext_RW0_addr ; 
             frontend_icache_tag_array_0_ext__RW0_ren_d0  <= frontend_icache_tag_array_0_ext_RW0_en ; 
             frontend_icache_tag_array_0_ext__RW0_rmode_d0  <= frontend_icache_tag_array_0_ext_RW0_wmode ;
             if ( frontend_icache_tag_array_0_ext_RW0_en & frontend_icache_tag_array_0_ext_RW0_wmode &1'h1) 
                 frontend_icache_tag_array_0_ext_Memory  [ frontend_icache_tag_array_0_ext_RW0_addr ]<= frontend_icache_tag_array_0_ext_RW0_wdata ;
         end
  assign  frontend_icache_tag_array_0_ext_RW0_rdata = frontend_icache_tag_array_0_ext__RW0_ren_d0 &~ frontend_icache_tag_array_0_ext__RW0_rmode_d0  ?  frontend_icache_tag_array_0_ext_Memory [ frontend_icache_tag_array_0_ext__RW0_raddr_d0 ]:21'bx;
    assign frontend_icache_tag_array_0_ext_RW0_addr = frontend_icache_refill_done ? frontend_icache_refill_idx:frontend_icache__tag_rdata_T_4;
    assign frontend_icache_tag_array_0_ext_RW0_en = frontend_icache_readEnable_0|frontend_icache_refill_done;
    assign frontend_icache_tag_array_0_ext_RW0_clk = frontend_icache_clock;
    assign frontend_icache_tag_array_0_ext_RW0_wmode = frontend_icache_refill_done;
    assign frontend_icache_tag_array_0_ext_RW0_wdata = frontend_icache_enc_tag;
    assign frontend_icache__tag_array_0_ext_RW0_rdata = frontend_icache_tag_array_0_ext_RW0_rdata;
      
    wire[9:0] frontend_icache_data_arrays_0_0_ext_RW0_addr;
    wire frontend_icache_data_arrays_0_0_ext_RW0_en;
    wire frontend_icache_data_arrays_0_0_ext_RW0_clk;
    wire frontend_icache_data_arrays_0_0_ext_RW0_wmode;
    wire[31:0] frontend_icache_data_arrays_0_0_ext_RW0_wdata;
    wire[31:0] frontend_icache_data_arrays_0_0_ext_RW0_rdata;

    reg[31:0] frontend_icache_data_arrays_0_0_ext_Memory [0:1023]; reg[9:0] frontend_icache_data_arrays_0_0_ext__RW0_raddr_d0 ; 
    reg frontend_icache_data_arrays_0_0_ext__RW0_ren_d0 ; 
    reg frontend_icache_data_arrays_0_0_ext__RW0_rmode_d0 ; 
  always @( posedge  frontend_icache_data_arrays_0_0_ext_RW0_clk )
         begin  
             frontend_icache_data_arrays_0_0_ext__RW0_raddr_d0  <= frontend_icache_data_arrays_0_0_ext_RW0_addr ; 
             frontend_icache_data_arrays_0_0_ext__RW0_ren_d0  <= frontend_icache_data_arrays_0_0_ext_RW0_en ; 
             frontend_icache_data_arrays_0_0_ext__RW0_rmode_d0  <= frontend_icache_data_arrays_0_0_ext_RW0_wmode ;
             if ( frontend_icache_data_arrays_0_0_ext_RW0_en & frontend_icache_data_arrays_0_0_ext_RW0_wmode &1'h1) 
                 frontend_icache_data_arrays_0_0_ext_Memory  [ frontend_icache_data_arrays_0_0_ext_RW0_addr ]<= frontend_icache_data_arrays_0_0_ext_RW0_wdata ;
         end
  assign  frontend_icache_data_arrays_0_0_ext_RW0_rdata = frontend_icache_data_arrays_0_0_ext__RW0_ren_d0 &~ frontend_icache_data_arrays_0_0_ext__RW0_rmode_d0  ?  frontend_icache_data_arrays_0_0_ext_Memory [ frontend_icache_data_arrays_0_0_ext__RW0_raddr_d0 ]:32'bx;
    assign frontend_icache_data_arrays_0_0_ext_RW0_addr = frontend_icache_mem_idx;
    assign frontend_icache_data_arrays_0_0_ext_RW0_en = frontend_icache_readEnable|frontend_icache_wen;
    assign frontend_icache_data_arrays_0_0_ext_RW0_clk = frontend_icache_clock;
    assign frontend_icache_data_arrays_0_0_ext_RW0_wmode = frontend_icache_wen;
    assign frontend_icache_data_arrays_0_0_ext_RW0_wdata = frontend_icache_data;
    assign frontend_icache_s1_dout_0 = frontend_icache_data_arrays_0_0_ext_RW0_rdata;
     
  assign  frontend_icache_auto_master_out_a_valid = frontend_icache_masterNodeOut_a_valid ; 
  assign  frontend_icache_auto_master_out_a_bits_address = frontend_icache_masterNodeOut_a_bits_address ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_readalloc = frontend_icache_masterNodeOut_a_bits_user_amba_prot_readalloc ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_writealloc = frontend_icache_masterNodeOut_a_bits_user_amba_prot_writealloc ; 
  assign  frontend_icache_io_resp_valid = frontend_icache_s2_valid & frontend_icache_s2_hit ; 
  assign  frontend_icache_io_resp_bits_data = frontend_icache_s2_dout_0 ; 
  assign  frontend_icache_io_resp_bits_ae = frontend_icache_s2_tl_error ;
    assign frontend_icache_clock = frontend_clock;
    assign frontend_icache_reset = frontend_reset;
    assign frontend_icache_auto_master_out_a_ready = frontend_auto_icache_master_out_a_ready;
    assign frontend_auto_icache_master_out_a_valid = frontend_icache_auto_master_out_a_valid;
    assign frontend_auto_icache_master_out_a_bits_address = frontend_icache_auto_master_out_a_bits_address;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_readalloc = frontend_icache_auto_master_out_a_bits_user_amba_prot_readalloc;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_writealloc = frontend_icache_auto_master_out_a_bits_user_amba_prot_writealloc;
    assign frontend_icache_auto_master_out_d_valid = frontend_auto_icache_master_out_d_valid;
    assign frontend_icache_auto_master_out_d_bits_opcode = frontend_auto_icache_master_out_d_bits_opcode;
    assign frontend_icache_auto_master_out_d_bits_param = frontend_auto_icache_master_out_d_bits_param;
    assign frontend_icache_auto_master_out_d_bits_size = frontend_auto_icache_master_out_d_bits_size;
    assign frontend_icache_auto_master_out_d_bits_sink = frontend_auto_icache_master_out_d_bits_sink;
    assign frontend_icache_auto_master_out_d_bits_denied = frontend_auto_icache_master_out_d_bits_denied;
    assign frontend_icache_auto_master_out_d_bits_data = frontend_auto_icache_master_out_d_bits_data;
    assign frontend_icache_auto_master_out_d_bits_corrupt = frontend_auto_icache_master_out_d_bits_corrupt;
    assign frontend_icache_io_req_valid = frontend_s0_valid;
    assign frontend_icache_io_req_bits_addr = frontend__io_cpu_npc_T_3;
    assign frontend_icache_io_s1_paddr = frontend__tlb_io_resp_paddr;
    assign frontend_icache_io_s2_vaddr = frontend_s2_pc;
    assign frontend_icache_io_s1_kill = frontend_s2_redirect|frontend_s2_replay;
    assign frontend_icache_io_s2_kill = frontend__icache_io_s2_kill_T_2;
    assign frontend_icache_io_s2_cacheable = frontend_s2_tlb_resp_cacheable;
    assign frontend__icache_io_resp_valid = frontend_icache_io_resp_valid;
    assign frontend__icache_io_resp_bits_data = frontend_icache_io_resp_bits_data;
    assign frontend__icache_io_resp_bits_ae = frontend_icache_io_resp_bits_ae;
    assign frontend_icache_io_invalidate = frontend_io_cpu_flush_icache;
      
    wire frontend_fq_clock;
    wire frontend_fq_reset;
    wire frontend_fq_io_enq_ready;
    wire frontend_fq_io_enq_valid;
    wire[1:0] frontend_fq_io_enq_bits_btb_cfiType;
    wire[1:0] frontend_fq_io_enq_bits_btb_mask;
    wire frontend_fq_io_enq_bits_btb_bridx;
    wire[31:0] frontend_fq_io_enq_bits_btb_target;
    wire frontend_fq_io_enq_bits_btb_entry;
    wire[7:0] frontend_fq_io_enq_bits_btb_bht_history;
    wire frontend_fq_io_enq_bits_btb_bht_value;
    wire[31:0] frontend_fq_io_enq_bits_pc;
    wire[31:0] frontend_fq_io_enq_bits_data;
    wire[1:0] frontend_fq_io_enq_bits_mask;
    wire frontend_fq_io_enq_bits_xcpt_pf_inst;
    wire frontend_fq_io_enq_bits_xcpt_ae_inst;
    wire frontend_fq_io_enq_bits_replay;
    wire frontend_fq_io_deq_ready;
    wire frontend_fq_io_deq_valid;
    wire[1:0] frontend_fq_io_deq_bits_btb_cfiType;
    wire frontend_fq_io_deq_bits_btb_taken;
    wire[1:0] frontend_fq_io_deq_bits_btb_mask;
    wire frontend_fq_io_deq_bits_btb_bridx;
    wire[31:0] frontend_fq_io_deq_bits_btb_target;
    wire frontend_fq_io_deq_bits_btb_entry;
    wire[7:0] frontend_fq_io_deq_bits_btb_bht_history;
    wire frontend_fq_io_deq_bits_btb_bht_value;
    wire[31:0] frontend_fq_io_deq_bits_pc;
    wire[31:0] frontend_fq_io_deq_bits_data;
    wire[1:0] frontend_fq_io_deq_bits_mask;
    wire frontend_fq_io_deq_bits_xcpt_pf_inst;
    wire frontend_fq_io_deq_bits_xcpt_gf_inst;
    wire frontend_fq_io_deq_bits_xcpt_ae_inst;
    wire frontend_fq_io_deq_bits_replay;
    wire[4:0] frontend_fq_io_mask;

    wire frontend_fq_wdata_3_btb_taken =1'h0; 
    reg frontend_fq_valid_0 ; 
    reg frontend_fq_valid_1 ; 
    reg frontend_fq_valid_2 ; 
    reg frontend_fq_valid_3 ; 
    reg frontend_fq_valid_4 ; reg[1:0] frontend_fq_elts_0_btb_cfiType ; 
    reg frontend_fq_elts_0_btb_taken ; reg[1:0] frontend_fq_elts_0_btb_mask ; 
    reg frontend_fq_elts_0_btb_bridx ; reg[31:0] frontend_fq_elts_0_btb_target ; 
    reg frontend_fq_elts_0_btb_entry ; reg[7:0] frontend_fq_elts_0_btb_bht_history ; 
    reg frontend_fq_elts_0_btb_bht_value ; reg[31:0] frontend_fq_elts_0_pc ; reg[31:0] frontend_fq_elts_0_data ; reg[1:0] frontend_fq_elts_0_mask ; 
    reg frontend_fq_elts_0_xcpt_pf_inst ; 
    reg frontend_fq_elts_0_xcpt_gf_inst ; 
    reg frontend_fq_elts_0_xcpt_ae_inst ; 
    reg frontend_fq_elts_0_replay ; reg[1:0] frontend_fq_elts_1_btb_cfiType ; 
    reg frontend_fq_elts_1_btb_taken ; reg[1:0] frontend_fq_elts_1_btb_mask ; 
    reg frontend_fq_elts_1_btb_bridx ; reg[31:0] frontend_fq_elts_1_btb_target ; 
    reg frontend_fq_elts_1_btb_entry ; reg[7:0] frontend_fq_elts_1_btb_bht_history ; 
    reg frontend_fq_elts_1_btb_bht_value ; reg[31:0] frontend_fq_elts_1_pc ; reg[31:0] frontend_fq_elts_1_data ; reg[1:0] frontend_fq_elts_1_mask ; 
    reg frontend_fq_elts_1_xcpt_pf_inst ; 
    reg frontend_fq_elts_1_xcpt_gf_inst ; 
    reg frontend_fq_elts_1_xcpt_ae_inst ; 
    reg frontend_fq_elts_1_replay ; reg[1:0] frontend_fq_elts_2_btb_cfiType ; 
    reg frontend_fq_elts_2_btb_taken ; reg[1:0] frontend_fq_elts_2_btb_mask ; 
    reg frontend_fq_elts_2_btb_bridx ; reg[31:0] frontend_fq_elts_2_btb_target ; 
    reg frontend_fq_elts_2_btb_entry ; reg[7:0] frontend_fq_elts_2_btb_bht_history ; 
    reg frontend_fq_elts_2_btb_bht_value ; reg[31:0] frontend_fq_elts_2_pc ; reg[31:0] frontend_fq_elts_2_data ; reg[1:0] frontend_fq_elts_2_mask ; 
    reg frontend_fq_elts_2_xcpt_pf_inst ; 
    reg frontend_fq_elts_2_xcpt_gf_inst ; 
    reg frontend_fq_elts_2_xcpt_ae_inst ; 
    reg frontend_fq_elts_2_replay ; reg[1:0] frontend_fq_elts_3_btb_cfiType ; 
    reg frontend_fq_elts_3_btb_taken ; reg[1:0] frontend_fq_elts_3_btb_mask ; 
    reg frontend_fq_elts_3_btb_bridx ; reg[31:0] frontend_fq_elts_3_btb_target ; 
    reg frontend_fq_elts_3_btb_entry ; reg[7:0] frontend_fq_elts_3_btb_bht_history ; 
    reg frontend_fq_elts_3_btb_bht_value ; reg[31:0] frontend_fq_elts_3_pc ; reg[31:0] frontend_fq_elts_3_data ; reg[1:0] frontend_fq_elts_3_mask ; 
    reg frontend_fq_elts_3_xcpt_pf_inst ; 
    reg frontend_fq_elts_3_xcpt_gf_inst ; 
    reg frontend_fq_elts_3_xcpt_ae_inst ; 
    reg frontend_fq_elts_3_replay ; reg[1:0] frontend_fq_elts_4_btb_cfiType ; reg[1:0] frontend_fq_elts_4_btb_mask ; 
    reg frontend_fq_elts_4_btb_bridx ; reg[31:0] frontend_fq_elts_4_btb_target ; 
    reg frontend_fq_elts_4_btb_entry ; reg[7:0] frontend_fq_elts_4_btb_bht_history ; 
    reg frontend_fq_elts_4_btb_bht_value ; reg[31:0] frontend_fq_elts_4_pc ; reg[31:0] frontend_fq_elts_4_data ; reg[1:0] frontend_fq_elts_4_mask ; 
    reg frontend_fq_elts_4_xcpt_pf_inst ; 
    reg frontend_fq_elts_4_xcpt_gf_inst ; 
    reg frontend_fq_elts_4_xcpt_ae_inst ; 
    reg frontend_fq_elts_4_replay ; 
    wire[1:0] frontend_fq_wdata_btb_cfiType = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_btb_taken = frontend_fq_valid_1 & frontend_fq_elts_1_btb_taken ; 
    wire[1:0] frontend_fq_wdata_btb_mask = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_btb_bridx = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[31:0] frontend_fq_wdata_btb_target = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_btb_entry = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_btb_bht_history = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_btb_bht_value = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[31:0] frontend_fq_wdata_pc = frontend_fq_valid_1  ?  frontend_fq_elts_1_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_data = frontend_fq_valid_1  ?  frontend_fq_elts_1_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_mask = frontend_fq_valid_1  ?  frontend_fq_elts_1_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_xcpt_pf_inst = frontend_fq_valid_1  ?  frontend_fq_elts_1_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_xcpt_gf_inst = frontend_fq_valid_1 & frontend_fq_elts_1_xcpt_gf_inst ; 
    wire frontend_fq_wdata_xcpt_ae_inst = frontend_fq_valid_1  ?  frontend_fq_elts_1_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_replay = frontend_fq_valid_1  ?  frontend_fq_elts_1_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq__valid_4_T_4 =~ frontend_fq_valid_4 & frontend_fq_io_enq_valid ; 
    wire frontend_fq_wen = frontend_fq_io_deq_ready  ?  frontend_fq_valid_1 | frontend_fq__valid_4_T_4 & frontend_fq_valid_0 : frontend_fq__valid_4_T_4 &~ frontend_fq_valid_0 ; 
    wire[1:0] frontend_fq_wdata_1_btb_cfiType = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_1_btb_taken = frontend_fq_valid_2 & frontend_fq_elts_2_btb_taken ; 
    wire[1:0] frontend_fq_wdata_1_btb_mask = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_1_btb_bridx = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[31:0] frontend_fq_wdata_1_btb_target = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_1_btb_entry = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_1_btb_bht_history = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_1_btb_bht_value = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[31:0] frontend_fq_wdata_1_pc = frontend_fq_valid_2  ?  frontend_fq_elts_2_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_1_data = frontend_fq_valid_2  ?  frontend_fq_elts_2_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_1_mask = frontend_fq_valid_2  ?  frontend_fq_elts_2_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_1_xcpt_pf_inst = frontend_fq_valid_2  ?  frontend_fq_elts_2_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_1_xcpt_gf_inst = frontend_fq_valid_2 & frontend_fq_elts_2_xcpt_gf_inst ; 
    wire frontend_fq_wdata_1_xcpt_ae_inst = frontend_fq_valid_2  ?  frontend_fq_elts_2_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_1_replay = frontend_fq_valid_2  ?  frontend_fq_elts_2_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq_wen_1 = frontend_fq_io_deq_ready  ?  frontend_fq_valid_2 | frontend_fq__valid_4_T_4 & frontend_fq_valid_1 : frontend_fq__valid_4_T_4 & frontend_fq_valid_0 &~ frontend_fq_valid_1 ; 
    wire[1:0] frontend_fq_wdata_2_btb_cfiType = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_2_btb_taken = frontend_fq_valid_3 & frontend_fq_elts_3_btb_taken ; 
    wire[1:0] frontend_fq_wdata_2_btb_mask = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_2_btb_bridx = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[31:0] frontend_fq_wdata_2_btb_target = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_2_btb_entry = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_2_btb_bht_history = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_2_btb_bht_value = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[31:0] frontend_fq_wdata_2_pc = frontend_fq_valid_3  ?  frontend_fq_elts_3_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_2_data = frontend_fq_valid_3  ?  frontend_fq_elts_3_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_2_mask = frontend_fq_valid_3  ?  frontend_fq_elts_3_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_2_xcpt_pf_inst = frontend_fq_valid_3  ?  frontend_fq_elts_3_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_2_xcpt_gf_inst = frontend_fq_valid_3 & frontend_fq_elts_3_xcpt_gf_inst ; 
    wire frontend_fq_wdata_2_xcpt_ae_inst = frontend_fq_valid_3  ?  frontend_fq_elts_3_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_2_replay = frontend_fq_valid_3  ?  frontend_fq_elts_3_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq_wen_2 = frontend_fq_io_deq_ready  ?  frontend_fq_valid_3 | frontend_fq__valid_4_T_4 & frontend_fq_valid_2 : frontend_fq__valid_4_T_4 & frontend_fq_valid_1 &~ frontend_fq_valid_2 ; 
    wire[1:0] frontend_fq_wdata_3_btb_cfiType = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire[1:0] frontend_fq_wdata_3_btb_mask = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_3_btb_bridx = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[31:0] frontend_fq_wdata_3_btb_target = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_3_btb_entry = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_3_btb_bht_history = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_3_btb_bht_value = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[31:0] frontend_fq_wdata_3_pc = frontend_fq_valid_4  ?  frontend_fq_elts_4_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_3_data = frontend_fq_valid_4  ?  frontend_fq_elts_4_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_3_mask = frontend_fq_valid_4  ?  frontend_fq_elts_4_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_3_xcpt_pf_inst = frontend_fq_valid_4  ?  frontend_fq_elts_4_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_3_xcpt_gf_inst = frontend_fq_valid_4 & frontend_fq_elts_4_xcpt_gf_inst ; 
    wire frontend_fq_wdata_3_xcpt_ae_inst = frontend_fq_valid_4  ?  frontend_fq_elts_4_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_3_replay = frontend_fq_valid_4  ?  frontend_fq_elts_4_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq_wen_3 = frontend_fq_io_deq_ready  ?  frontend_fq_valid_4 | frontend_fq__valid_4_T_4 & frontend_fq_valid_3 : frontend_fq__valid_4_T_4 & frontend_fq_valid_2 &~ frontend_fq_valid_3 ; 
    wire frontend_fq_wen_4 = frontend_fq_io_deq_ready  ?  frontend_fq__valid_4_T_4 & frontend_fq_valid_4 : frontend_fq__valid_4_T_4 & frontend_fq_valid_3 &~ frontend_fq_valid_4 ; 
    wire[1:0] frontend_fq_io_mask_lo ={ frontend_fq_valid_1 , frontend_fq_valid_0 }; 
    wire[1:0] frontend_fq_io_mask_hi_hi ={ frontend_fq_valid_4 , frontend_fq_valid_3 }; 
    wire[2:0] frontend_fq_io_mask_hi ={ frontend_fq_io_mask_hi_hi , frontend_fq_valid_2 }; 
  always @( posedge  frontend_fq_clock )
         begin 
             if ( frontend_fq_reset )
                 begin  
                     frontend_fq_valid_0  <=1'h0; 
                     frontend_fq_valid_1  <=1'h0; 
                     frontend_fq_valid_2  <=1'h0; 
                     frontend_fq_valid_3  <=1'h0; 
                     frontend_fq_valid_4  <=1'h0;
                 end 
              else 
                 if ( frontend_fq_io_deq_ready )
                     begin  
                         frontend_fq_valid_0  <= frontend_fq_valid_1 | frontend_fq__valid_4_T_4 & frontend_fq_valid_0 ; 
                         frontend_fq_valid_1  <= frontend_fq_valid_2 | frontend_fq__valid_4_T_4 & frontend_fq_valid_1 ; 
                         frontend_fq_valid_2  <= frontend_fq_valid_3 | frontend_fq__valid_4_T_4 & frontend_fq_valid_2 ; 
                         frontend_fq_valid_3  <= frontend_fq_valid_4 | frontend_fq__valid_4_T_4 & frontend_fq_valid_3 ; 
                         frontend_fq_valid_4  <= frontend_fq__valid_4_T_4 & frontend_fq_valid_4 ;
                     end 
                  else 
                     begin  
                         frontend_fq_valid_0  <= frontend_fq__valid_4_T_4 | frontend_fq_valid_0 ; 
                         frontend_fq_valid_1  <= frontend_fq__valid_4_T_4 & frontend_fq_valid_0 | frontend_fq_valid_1 ; 
                         frontend_fq_valid_2  <= frontend_fq__valid_4_T_4 & frontend_fq_valid_1 | frontend_fq_valid_2 ; 
                         frontend_fq_valid_3  <= frontend_fq__valid_4_T_4 & frontend_fq_valid_2 | frontend_fq_valid_3 ; 
                         frontend_fq_valid_4  <= frontend_fq__valid_4_T_4 & frontend_fq_valid_3 | frontend_fq_valid_4 ;
                     end 
             if ( frontend_fq_wen )
                 begin  
                     frontend_fq_elts_0_btb_cfiType  <= frontend_fq_wdata_btb_cfiType ; 
                     frontend_fq_elts_0_btb_taken  <= frontend_fq_wdata_btb_taken ; 
                     frontend_fq_elts_0_btb_mask  <= frontend_fq_wdata_btb_mask ; 
                     frontend_fq_elts_0_btb_bridx  <= frontend_fq_wdata_btb_bridx ; 
                     frontend_fq_elts_0_btb_target  <= frontend_fq_wdata_btb_target ; 
                     frontend_fq_elts_0_btb_entry  <= frontend_fq_wdata_btb_entry ; 
                     frontend_fq_elts_0_btb_bht_history  <= frontend_fq_wdata_btb_bht_history ; 
                     frontend_fq_elts_0_btb_bht_value  <= frontend_fq_wdata_btb_bht_value ; 
                     frontend_fq_elts_0_pc  <= frontend_fq_wdata_pc ; 
                     frontend_fq_elts_0_data  <= frontend_fq_wdata_data ; 
                     frontend_fq_elts_0_mask  <= frontend_fq_wdata_mask ; 
                     frontend_fq_elts_0_xcpt_pf_inst  <= frontend_fq_wdata_xcpt_pf_inst ; 
                     frontend_fq_elts_0_xcpt_gf_inst  <= frontend_fq_wdata_xcpt_gf_inst ; 
                     frontend_fq_elts_0_xcpt_ae_inst  <= frontend_fq_wdata_xcpt_ae_inst ; 
                     frontend_fq_elts_0_replay  <= frontend_fq_wdata_replay ;
                 end 
             if ( frontend_fq_wen_1 )
                 begin  
                     frontend_fq_elts_1_btb_cfiType  <= frontend_fq_wdata_1_btb_cfiType ; 
                     frontend_fq_elts_1_btb_taken  <= frontend_fq_wdata_1_btb_taken ; 
                     frontend_fq_elts_1_btb_mask  <= frontend_fq_wdata_1_btb_mask ; 
                     frontend_fq_elts_1_btb_bridx  <= frontend_fq_wdata_1_btb_bridx ; 
                     frontend_fq_elts_1_btb_target  <= frontend_fq_wdata_1_btb_target ; 
                     frontend_fq_elts_1_btb_entry  <= frontend_fq_wdata_1_btb_entry ; 
                     frontend_fq_elts_1_btb_bht_history  <= frontend_fq_wdata_1_btb_bht_history ; 
                     frontend_fq_elts_1_btb_bht_value  <= frontend_fq_wdata_1_btb_bht_value ; 
                     frontend_fq_elts_1_pc  <= frontend_fq_wdata_1_pc ; 
                     frontend_fq_elts_1_data  <= frontend_fq_wdata_1_data ; 
                     frontend_fq_elts_1_mask  <= frontend_fq_wdata_1_mask ; 
                     frontend_fq_elts_1_xcpt_pf_inst  <= frontend_fq_wdata_1_xcpt_pf_inst ; 
                     frontend_fq_elts_1_xcpt_gf_inst  <= frontend_fq_wdata_1_xcpt_gf_inst ; 
                     frontend_fq_elts_1_xcpt_ae_inst  <= frontend_fq_wdata_1_xcpt_ae_inst ; 
                     frontend_fq_elts_1_replay  <= frontend_fq_wdata_1_replay ;
                 end 
             if ( frontend_fq_wen_2 )
                 begin  
                     frontend_fq_elts_2_btb_cfiType  <= frontend_fq_wdata_2_btb_cfiType ; 
                     frontend_fq_elts_2_btb_taken  <= frontend_fq_wdata_2_btb_taken ; 
                     frontend_fq_elts_2_btb_mask  <= frontend_fq_wdata_2_btb_mask ; 
                     frontend_fq_elts_2_btb_bridx  <= frontend_fq_wdata_2_btb_bridx ; 
                     frontend_fq_elts_2_btb_target  <= frontend_fq_wdata_2_btb_target ; 
                     frontend_fq_elts_2_btb_entry  <= frontend_fq_wdata_2_btb_entry ; 
                     frontend_fq_elts_2_btb_bht_history  <= frontend_fq_wdata_2_btb_bht_history ; 
                     frontend_fq_elts_2_btb_bht_value  <= frontend_fq_wdata_2_btb_bht_value ; 
                     frontend_fq_elts_2_pc  <= frontend_fq_wdata_2_pc ; 
                     frontend_fq_elts_2_data  <= frontend_fq_wdata_2_data ; 
                     frontend_fq_elts_2_mask  <= frontend_fq_wdata_2_mask ; 
                     frontend_fq_elts_2_xcpt_pf_inst  <= frontend_fq_wdata_2_xcpt_pf_inst ; 
                     frontend_fq_elts_2_xcpt_gf_inst  <= frontend_fq_wdata_2_xcpt_gf_inst ; 
                     frontend_fq_elts_2_xcpt_ae_inst  <= frontend_fq_wdata_2_xcpt_ae_inst ; 
                     frontend_fq_elts_2_replay  <= frontend_fq_wdata_2_replay ;
                 end 
             if ( frontend_fq_wen_3 )
                 begin  
                     frontend_fq_elts_3_btb_cfiType  <= frontend_fq_wdata_3_btb_cfiType ; 
                     frontend_fq_elts_3_btb_mask  <= frontend_fq_wdata_3_btb_mask ; 
                     frontend_fq_elts_3_btb_bridx  <= frontend_fq_wdata_3_btb_bridx ; 
                     frontend_fq_elts_3_btb_target  <= frontend_fq_wdata_3_btb_target ; 
                     frontend_fq_elts_3_btb_entry  <= frontend_fq_wdata_3_btb_entry ; 
                     frontend_fq_elts_3_btb_bht_history  <= frontend_fq_wdata_3_btb_bht_history ; 
                     frontend_fq_elts_3_btb_bht_value  <= frontend_fq_wdata_3_btb_bht_value ; 
                     frontend_fq_elts_3_pc  <= frontend_fq_wdata_3_pc ; 
                     frontend_fq_elts_3_data  <= frontend_fq_wdata_3_data ; 
                     frontend_fq_elts_3_mask  <= frontend_fq_wdata_3_mask ; 
                     frontend_fq_elts_3_xcpt_pf_inst  <= frontend_fq_wdata_3_xcpt_pf_inst ; 
                     frontend_fq_elts_3_xcpt_gf_inst  <= frontend_fq_wdata_3_xcpt_gf_inst ; 
                     frontend_fq_elts_3_xcpt_ae_inst  <= frontend_fq_wdata_3_xcpt_ae_inst ; 
                     frontend_fq_elts_3_replay  <= frontend_fq_wdata_3_replay ;
                 end  
             frontend_fq_elts_3_btb_taken  <=~ frontend_fq_wen_3 & frontend_fq_elts_3_btb_taken ;
             if ( frontend_fq_wen_4 )
                 begin  
                     frontend_fq_elts_4_btb_cfiType  <= frontend_fq_io_enq_bits_btb_cfiType ; 
                     frontend_fq_elts_4_btb_mask  <= frontend_fq_io_enq_bits_btb_mask ; 
                     frontend_fq_elts_4_btb_bridx  <= frontend_fq_io_enq_bits_btb_bridx ; 
                     frontend_fq_elts_4_btb_target  <= frontend_fq_io_enq_bits_btb_target ; 
                     frontend_fq_elts_4_btb_entry  <= frontend_fq_io_enq_bits_btb_entry ; 
                     frontend_fq_elts_4_btb_bht_history  <= frontend_fq_io_enq_bits_btb_bht_history ; 
                     frontend_fq_elts_4_btb_bht_value  <= frontend_fq_io_enq_bits_btb_bht_value ; 
                     frontend_fq_elts_4_pc  <= frontend_fq_io_enq_bits_pc ; 
                     frontend_fq_elts_4_data  <= frontend_fq_io_enq_bits_data ; 
                     frontend_fq_elts_4_mask  <= frontend_fq_io_enq_bits_mask ; 
                     frontend_fq_elts_4_xcpt_pf_inst  <= frontend_fq_io_enq_bits_xcpt_pf_inst ; 
                     frontend_fq_elts_4_xcpt_ae_inst  <= frontend_fq_io_enq_bits_xcpt_ae_inst ; 
                     frontend_fq_elts_4_replay  <= frontend_fq_io_enq_bits_replay ;
                 end  
             frontend_fq_elts_4_xcpt_gf_inst  <=~ frontend_fq_wen_4 & frontend_fq_elts_4_xcpt_gf_inst ;
         end
  assign  frontend_fq_io_enq_ready =~ frontend_fq_valid_4 ; 
  assign  frontend_fq_io_deq_valid = frontend_fq_io_enq_valid | frontend_fq_valid_0 ; 
  assign  frontend_fq_io_deq_bits_btb_cfiType = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
  assign  frontend_fq_io_deq_bits_btb_taken = frontend_fq_valid_0 & frontend_fq_elts_0_btb_taken ; 
  assign  frontend_fq_io_deq_bits_btb_mask = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
  assign  frontend_fq_io_deq_bits_btb_bridx = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
  assign  frontend_fq_io_deq_bits_btb_target = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_target : frontend_fq_io_enq_bits_btb_target ; 
  assign  frontend_fq_io_deq_bits_btb_entry = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
  assign  frontend_fq_io_deq_bits_btb_bht_history = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
  assign  frontend_fq_io_deq_bits_btb_bht_value = frontend_fq_valid_0  ?  frontend_fq_elts_0_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
  assign  frontend_fq_io_deq_bits_pc = frontend_fq_valid_0  ?  frontend_fq_elts_0_pc : frontend_fq_io_enq_bits_pc ; 
  assign  frontend_fq_io_deq_bits_data = frontend_fq_valid_0  ?  frontend_fq_elts_0_data : frontend_fq_io_enq_bits_data ; 
  assign  frontend_fq_io_deq_bits_mask = frontend_fq_valid_0  ?  frontend_fq_elts_0_mask : frontend_fq_io_enq_bits_mask ; 
  assign  frontend_fq_io_deq_bits_xcpt_pf_inst = frontend_fq_valid_0  ?  frontend_fq_elts_0_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
  assign  frontend_fq_io_deq_bits_xcpt_gf_inst = frontend_fq_valid_0 & frontend_fq_elts_0_xcpt_gf_inst ; 
  assign  frontend_fq_io_deq_bits_xcpt_ae_inst = frontend_fq_valid_0  ?  frontend_fq_elts_0_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
  assign  frontend_fq_io_deq_bits_replay = frontend_fq_valid_0  ?  frontend_fq_elts_0_replay : frontend_fq_io_enq_bits_replay ; 
  assign  frontend_fq_io_mask ={ frontend_fq_io_mask_hi , frontend_fq_io_mask_lo };
    assign frontend_fq_clock = frontend_clock;
    assign frontend_fq_reset = frontend_reset|frontend_io_cpu_req_valid;
    assign frontend__fq_io_enq_ready = frontend_fq_io_enq_ready;
    assign frontend_fq_io_enq_valid = frontend__fq_io_enq_valid_T_6;
    assign frontend_fq_io_enq_bits_btb_cfiType = 2'h0;
    assign frontend_fq_io_enq_bits_btb_mask = 2'h0;
    assign frontend_fq_io_enq_bits_btb_bridx = 1'h0;
    assign frontend_fq_io_enq_bits_btb_target = 32'h0;
    assign frontend_fq_io_enq_bits_btb_entry = 1'h0;
    assign frontend_fq_io_enq_bits_btb_bht_history = 8'h0;
    assign frontend_fq_io_enq_bits_btb_bht_value = 1'h0;
    assign frontend_fq_io_enq_bits_pc = frontend_s2_pc;
    assign frontend_fq_io_enq_bits_data = frontend__icache_io_resp_bits_data;
    assign frontend_fq_io_enq_bits_mask = frontend__fq_io_enq_bits_mask_T_1[1:0];
    assign frontend_fq_io_enq_bits_xcpt_pf_inst = frontend_s2_tlb_resp_pf_inst;
    assign frontend_fq_io_enq_bits_xcpt_ae_inst = frontend__icache_io_resp_valid&frontend__icache_io_resp_bits_ae|frontend_s2_tlb_resp_ae_inst;
    assign frontend_fq_io_enq_bits_replay = frontend__icache_io_s2_kill_T_2&~frontend__icache_io_resp_valid&~frontend_s2_xcpt;
    assign frontend_fq_io_deq_ready = frontend_io_cpu_resp_ready;
    assign frontend_io_cpu_resp_valid = frontend_fq_io_deq_valid;
    assign frontend_io_cpu_resp_bits_btb_cfiType = frontend_fq_io_deq_bits_btb_cfiType;
    assign frontend_io_cpu_resp_bits_btb_taken = frontend_fq_io_deq_bits_btb_taken;
    assign frontend_io_cpu_resp_bits_btb_mask = frontend_fq_io_deq_bits_btb_mask;
    assign frontend_io_cpu_resp_bits_btb_bridx = frontend_fq_io_deq_bits_btb_bridx;
    assign frontend_io_cpu_resp_bits_btb_target = frontend_fq_io_deq_bits_btb_target;
    assign frontend_io_cpu_resp_bits_btb_entry = frontend_fq_io_deq_bits_btb_entry;
    assign frontend_io_cpu_resp_bits_btb_bht_history = frontend_fq_io_deq_bits_btb_bht_history;
    assign frontend_io_cpu_resp_bits_btb_bht_value = frontend_fq_io_deq_bits_btb_bht_value;
    assign frontend_io_cpu_resp_bits_pc = frontend_fq_io_deq_bits_pc;
    assign frontend_io_cpu_resp_bits_data = frontend_fq_io_deq_bits_data;
    assign frontend_io_cpu_resp_bits_mask = frontend_fq_io_deq_bits_mask;
    assign frontend_io_cpu_resp_bits_xcpt_pf_inst = frontend_fq_io_deq_bits_xcpt_pf_inst;
    assign frontend_io_cpu_resp_bits_xcpt_gf_inst = frontend_fq_io_deq_bits_xcpt_gf_inst;
    assign frontend_io_cpu_resp_bits_xcpt_ae_inst = frontend_fq_io_deq_bits_xcpt_ae_inst;
    assign frontend_io_cpu_resp_bits_replay = frontend_fq_io_deq_bits_replay;
    assign frontend__fq_io_mask = frontend_fq_io_mask;
      
    wire[31:0] frontend_tlb_io_req_bits_vaddr;
    wire[31:0] frontend_tlb_io_resp_paddr;
    wire[31:0] frontend_tlb_io_resp_gpa;
    wire frontend_tlb_io_resp_pf_ld;
    wire frontend_tlb_io_resp_pf_inst;
    wire frontend_tlb_io_resp_ae_ld;
    wire frontend_tlb_io_resp_ae_inst;
    wire frontend_tlb_io_resp_ma_ld;
    wire frontend_tlb_io_resp_cacheable;
    wire frontend_tlb_io_resp_prefetchable;
    wire frontend_tlb_io_sfence_valid;
    wire frontend_tlb_io_ptw_req_bits_valid;
    wire[19:0] frontend_tlb_io_ptw_req_bits_bits_addr;
    wire frontend_tlb_io_ptw_req_bits_bits_need_gpa;
    wire frontend_tlb_io_ptw_req_bits_bits_vstage1;
    wire frontend_tlb_io_ptw_req_bits_bits_stage2;
    wire frontend_tlb_io_ptw_resp_bits_ae_ptw;
    wire frontend_tlb_io_ptw_resp_bits_ae_final;
    wire frontend_tlb_io_ptw_resp_bits_pf;
    wire frontend_tlb_io_ptw_resp_bits_gf;
    wire frontend_tlb_io_ptw_resp_bits_hr;
    wire frontend_tlb_io_ptw_resp_bits_hw;
    wire frontend_tlb_io_ptw_resp_bits_hx;
    wire[43:0] frontend_tlb_io_ptw_resp_bits_pte_ppn;
    wire frontend_tlb_io_ptw_resp_bits_pte_d;
    wire frontend_tlb_io_ptw_resp_bits_pte_a;
    wire frontend_tlb_io_ptw_resp_bits_pte_g;
    wire frontend_tlb_io_ptw_resp_bits_pte_u;
    wire frontend_tlb_io_ptw_resp_bits_pte_x;
    wire frontend_tlb_io_ptw_resp_bits_pte_w;
    wire frontend_tlb_io_ptw_resp_bits_pte_r;
    wire frontend_tlb_io_ptw_resp_bits_pte_v;
    wire frontend_tlb_io_ptw_resp_bits_gpa_is_pte;
    wire frontend_tlb_io_ptw_status_debug;
    wire frontend_tlb_io_ptw_pmp_0_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_0_cfg_a;
    wire frontend_tlb_io_ptw_pmp_0_cfg_x;
    wire frontend_tlb_io_ptw_pmp_0_cfg_w;
    wire frontend_tlb_io_ptw_pmp_0_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_0_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_0_mask;
    wire frontend_tlb_io_ptw_pmp_1_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_1_cfg_a;
    wire frontend_tlb_io_ptw_pmp_1_cfg_x;
    wire frontend_tlb_io_ptw_pmp_1_cfg_w;
    wire frontend_tlb_io_ptw_pmp_1_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_1_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_1_mask;
    wire frontend_tlb_io_ptw_pmp_2_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_2_cfg_a;
    wire frontend_tlb_io_ptw_pmp_2_cfg_x;
    wire frontend_tlb_io_ptw_pmp_2_cfg_w;
    wire frontend_tlb_io_ptw_pmp_2_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_2_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_2_mask;
    wire frontend_tlb_io_ptw_pmp_3_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_3_cfg_a;
    wire frontend_tlb_io_ptw_pmp_3_cfg_x;
    wire frontend_tlb_io_ptw_pmp_3_cfg_w;
    wire frontend_tlb_io_ptw_pmp_3_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_3_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_3_mask;
    wire frontend_tlb_io_ptw_pmp_4_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_4_cfg_a;
    wire frontend_tlb_io_ptw_pmp_4_cfg_x;
    wire frontend_tlb_io_ptw_pmp_4_cfg_w;
    wire frontend_tlb_io_ptw_pmp_4_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_4_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_4_mask;
    wire frontend_tlb_io_ptw_pmp_5_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_5_cfg_a;
    wire frontend_tlb_io_ptw_pmp_5_cfg_x;
    wire frontend_tlb_io_ptw_pmp_5_cfg_w;
    wire frontend_tlb_io_ptw_pmp_5_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_5_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_5_mask;
    wire frontend_tlb_io_ptw_pmp_6_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_6_cfg_a;
    wire frontend_tlb_io_ptw_pmp_6_cfg_x;
    wire frontend_tlb_io_ptw_pmp_6_cfg_w;
    wire frontend_tlb_io_ptw_pmp_6_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_6_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_6_mask;
    wire frontend_tlb_io_ptw_pmp_7_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_7_cfg_a;
    wire frontend_tlb_io_ptw_pmp_7_cfg_x;
    wire frontend_tlb_io_ptw_pmp_7_cfg_w;
    wire frontend_tlb_io_ptw_pmp_7_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_7_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_7_mask;
    wire frontend_tlb_io_kill;

    wire frontend_tlb__entries_barrier_5_io_y_u ; 
    wire frontend_tlb__entries_barrier_5_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_5_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_5_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_5_io_y_pf ; 
    wire frontend_tlb__entries_barrier_5_io_y_gf ; 
    wire frontend_tlb__entries_barrier_5_io_y_sw ; 
    wire frontend_tlb__entries_barrier_5_io_y_sx ; 
    wire frontend_tlb__entries_barrier_5_io_y_sr ; 
    wire frontend_tlb__entries_barrier_5_io_y_hw ; 
    wire frontend_tlb__entries_barrier_5_io_y_hx ; 
    wire frontend_tlb__entries_barrier_5_io_y_hr ; 
    wire frontend_tlb__entries_barrier_4_io_y_u ; 
    wire frontend_tlb__entries_barrier_4_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_4_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_4_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_4_io_y_pf ; 
    wire frontend_tlb__entries_barrier_4_io_y_gf ; 
    wire frontend_tlb__entries_barrier_4_io_y_sw ; 
    wire frontend_tlb__entries_barrier_4_io_y_sx ; 
    wire frontend_tlb__entries_barrier_4_io_y_sr ; 
    wire frontend_tlb__entries_barrier_4_io_y_hw ; 
    wire frontend_tlb__entries_barrier_4_io_y_hx ; 
    wire frontend_tlb__entries_barrier_4_io_y_hr ; 
    wire frontend_tlb__entries_barrier_4_io_y_pw ; 
    wire frontend_tlb__entries_barrier_4_io_y_px ; 
    wire frontend_tlb__entries_barrier_4_io_y_pr ; 
    wire frontend_tlb__entries_barrier_4_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_4_io_y_pal ; 
    wire frontend_tlb__entries_barrier_4_io_y_paa ; 
    wire frontend_tlb__entries_barrier_4_io_y_eff ; 
    wire frontend_tlb__entries_barrier_4_io_y_c ; 
    wire frontend_tlb__entries_barrier_3_io_y_u ; 
    wire frontend_tlb__entries_barrier_3_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_3_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_3_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_3_io_y_pf ; 
    wire frontend_tlb__entries_barrier_3_io_y_gf ; 
    wire frontend_tlb__entries_barrier_3_io_y_sw ; 
    wire frontend_tlb__entries_barrier_3_io_y_sx ; 
    wire frontend_tlb__entries_barrier_3_io_y_sr ; 
    wire frontend_tlb__entries_barrier_3_io_y_hw ; 
    wire frontend_tlb__entries_barrier_3_io_y_hx ; 
    wire frontend_tlb__entries_barrier_3_io_y_hr ; 
    wire frontend_tlb__entries_barrier_3_io_y_pw ; 
    wire frontend_tlb__entries_barrier_3_io_y_px ; 
    wire frontend_tlb__entries_barrier_3_io_y_pr ; 
    wire frontend_tlb__entries_barrier_3_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_3_io_y_pal ; 
    wire frontend_tlb__entries_barrier_3_io_y_paa ; 
    wire frontend_tlb__entries_barrier_3_io_y_eff ; 
    wire frontend_tlb__entries_barrier_3_io_y_c ; 
    wire frontend_tlb__entries_barrier_2_io_y_u ; 
    wire frontend_tlb__entries_barrier_2_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_2_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_2_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_2_io_y_pf ; 
    wire frontend_tlb__entries_barrier_2_io_y_gf ; 
    wire frontend_tlb__entries_barrier_2_io_y_sw ; 
    wire frontend_tlb__entries_barrier_2_io_y_sx ; 
    wire frontend_tlb__entries_barrier_2_io_y_sr ; 
    wire frontend_tlb__entries_barrier_2_io_y_hw ; 
    wire frontend_tlb__entries_barrier_2_io_y_hx ; 
    wire frontend_tlb__entries_barrier_2_io_y_hr ; 
    wire frontend_tlb__entries_barrier_2_io_y_pw ; 
    wire frontend_tlb__entries_barrier_2_io_y_px ; 
    wire frontend_tlb__entries_barrier_2_io_y_pr ; 
    wire frontend_tlb__entries_barrier_2_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_2_io_y_pal ; 
    wire frontend_tlb__entries_barrier_2_io_y_paa ; 
    wire frontend_tlb__entries_barrier_2_io_y_eff ; 
    wire frontend_tlb__entries_barrier_2_io_y_c ; 
    wire frontend_tlb__entries_barrier_1_io_y_u ; 
    wire frontend_tlb__entries_barrier_1_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_1_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_1_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_1_io_y_pf ; 
    wire frontend_tlb__entries_barrier_1_io_y_gf ; 
    wire frontend_tlb__entries_barrier_1_io_y_sw ; 
    wire frontend_tlb__entries_barrier_1_io_y_sx ; 
    wire frontend_tlb__entries_barrier_1_io_y_sr ; 
    wire frontend_tlb__entries_barrier_1_io_y_hw ; 
    wire frontend_tlb__entries_barrier_1_io_y_hx ; 
    wire frontend_tlb__entries_barrier_1_io_y_hr ; 
    wire frontend_tlb__entries_barrier_1_io_y_pw ; 
    wire frontend_tlb__entries_barrier_1_io_y_px ; 
    wire frontend_tlb__entries_barrier_1_io_y_pr ; 
    wire frontend_tlb__entries_barrier_1_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_1_io_y_pal ; 
    wire frontend_tlb__entries_barrier_1_io_y_paa ; 
    wire frontend_tlb__entries_barrier_1_io_y_eff ; 
    wire frontend_tlb__entries_barrier_1_io_y_c ; 
    wire frontend_tlb__entries_barrier_io_y_u ; 
    wire frontend_tlb__entries_barrier_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_io_y_pf ; 
    wire frontend_tlb__entries_barrier_io_y_gf ; 
    wire frontend_tlb__entries_barrier_io_y_sw ; 
    wire frontend_tlb__entries_barrier_io_y_sx ; 
    wire frontend_tlb__entries_barrier_io_y_sr ; 
    wire frontend_tlb__entries_barrier_io_y_hw ; 
    wire frontend_tlb__entries_barrier_io_y_hx ; 
    wire frontend_tlb__entries_barrier_io_y_hr ; 
    wire frontend_tlb__entries_barrier_io_y_pw ; 
    wire frontend_tlb__entries_barrier_io_y_px ; 
    wire frontend_tlb__entries_barrier_io_y_pr ; 
    wire frontend_tlb__entries_barrier_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_io_y_pal ; 
    wire frontend_tlb__entries_barrier_io_y_paa ; 
    wire frontend_tlb__entries_barrier_io_y_eff ; 
    wire frontend_tlb__entries_barrier_io_y_c ; 
    wire frontend_tlb__pmp_io_r ; 
    wire frontend_tlb__pmp_io_w ; 
    wire frontend_tlb__pmp_io_x ; 
    wire frontend_tlb_invalidate_refill = frontend_tlb_io_sfence_valid ; 
    wire frontend_tlb_newEntry_u = frontend_tlb_io_ptw_resp_bits_pte_u ; 
    wire frontend_tlb_newEntry_ae_ptw = frontend_tlb_io_ptw_resp_bits_ae_ptw ; 
    wire frontend_tlb_newEntry_ae_final = frontend_tlb_io_ptw_resp_bits_ae_final ; 
    wire frontend_tlb_newEntry_pf = frontend_tlb_io_ptw_resp_bits_pf ; 
    wire frontend_tlb_newEntry_gf = frontend_tlb_io_ptw_resp_bits_gf ; 
    wire frontend_tlb_newEntry_hw = frontend_tlb_io_ptw_resp_bits_hw ; 
    wire frontend_tlb_newEntry_hx = frontend_tlb_io_ptw_resp_bits_hx ; 
    wire frontend_tlb_newEntry_hr = frontend_tlb_io_ptw_resp_bits_hr ; 
    wire frontend_tlb_priv_s =1'h1; 
    wire frontend_tlb_cmd_read =1'h1; 
    wire[5:0] frontend_tlb_real_hits =6'h0; 
    wire[5:0] frontend_tlb_stage1_bypass =6'h0; 
    wire frontend_tlb_priv_v =1'h0; 
    wire frontend_tlb_priv_uses_vm =1'h0; 
    wire frontend_tlb_satp_mode =1'h0; 
    wire frontend_tlb_stage1_en =1'h0; 
    wire frontend_tlb_vstage1_en =1'h0; 
    wire frontend_tlb_stage2_en =1'h0; 
    wire frontend_tlb_vm_enabled =1'h0; 
    wire frontend_tlb_vsatp_mode_mismatch =1'h0; 
    wire frontend_tlb_do_refill =1'h0; 
    wire frontend_tlb_cacheable =1'h0; 
    wire frontend_tlb_sector_hits_0 =1'h0; 
    wire frontend_tlb_superpage_hits_0 =1'h0; 
    wire frontend_tlb_superpage_hits_1 =1'h0; 
    wire frontend_tlb_superpage_hits_2 =1'h0; 
    wire frontend_tlb_superpage_hits_3 =1'h0; 
    wire frontend_tlb_hitsVec_0 =1'h0; 
    wire frontend_tlb_hitsVec_1 =1'h0; 
    wire frontend_tlb_hitsVec_2 =1'h0; 
    wire frontend_tlb_hitsVec_3 =1'h0; 
    wire frontend_tlb_hitsVec_4 =1'h0; 
    wire frontend_tlb_hitsVec_5 =1'h0; 
    wire frontend_tlb_refill_v =1'h0; 
    wire frontend_tlb_newEntry_ae_stage2 =1'h0; 
    wire frontend_tlb_newEntry_c =1'h0; 
    wire frontend_tlb_newEntry_fragmented_superpage =1'h0; 
    wire frontend_tlb_sum =1'h0; 
    wire frontend_tlb_mxr =1'h0; 
    wire frontend_tlb_cmd_lrsc =1'h0; 
    wire frontend_tlb_cmd_amo_logical =1'h0; 
    wire frontend_tlb_cmd_amo_arithmetic =1'h0; 
    wire frontend_tlb_cmd_put_partial =1'h0; 
    wire frontend_tlb_cmd_readx =1'h0; 
    wire frontend_tlb_cmd_write =1'h0; 
    wire frontend_tlb_cmd_write_perms =1'h0; 
    wire frontend_tlb_tlb_hit_if_not_gpa_miss =1'h0; 
    wire frontend_tlb_tlb_hit =1'h0; 
    wire frontend_tlb_tlb_miss =1'h0; 
    wire frontend_tlb_state_reg_left_subtree_state =1'h0; 
    wire frontend_tlb_state_reg_right_subtree_state =1'h0; 
    wire frontend_tlb_multipleHits_leftOne =1'h0; 
    wire frontend_tlb_multipleHits_leftOne_1 =1'h0; 
    wire frontend_tlb_multipleHits_rightOne =1'h0; 
    wire frontend_tlb_multipleHits_rightOne_1 =1'h0; 
    wire frontend_tlb_multipleHits_rightTwo =1'h0; 
    wire frontend_tlb_multipleHits_leftOne_2 =1'h0; 
    wire frontend_tlb_multipleHits_leftTwo =1'h0; 
    wire frontend_tlb_multipleHits_leftOne_3 =1'h0; 
    wire frontend_tlb_multipleHits_leftOne_4 =1'h0; 
    wire frontend_tlb_multipleHits_rightOne_2 =1'h0; 
    wire frontend_tlb_multipleHits_rightOne_3 =1'h0; 
    wire frontend_tlb_multipleHits_rightTwo_1 =1'h0; 
    wire frontend_tlb_multipleHits_rightOne_4 =1'h0; 
    wire frontend_tlb_multipleHits_rightTwo_2 =1'h0; 
    wire frontend_tlb_multipleHits =1'h0; 
    wire[1:0] frontend_tlb_real_hits_lo_hi =2'h0; 
    wire[1:0] frontend_tlb_real_hits_hi_hi =2'h0; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_lo_lo =2'h0; 
    wire[1:0] frontend_tlb_waddr =2'h0; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_lo_lo =2'h0; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_lo_lo =2'h0; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_lo_lo =2'h0; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_lo_lo =2'h0; 
    wire[1:0] frontend_tlb_idx =2'h0; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_lo_lo =2'h0; 
    wire[2:0] frontend_tlb_real_hits_lo =3'h0; 
    wire[2:0] frontend_tlb_real_hits_hi =3'h0; 
    wire[6:0] frontend_tlb_hits =7'h40; 
    wire[6:0] frontend_tlb_hr_array =7'h7F; 
    wire[6:0] frontend_tlb_hw_array =7'h7F; 
    wire[6:0] frontend_tlb_hx_array =7'h7F; 
    wire[6:0] frontend_tlb_lrscAllowed =7'h0; 
    wire[6:0] frontend_tlb_ae_st_array =7'h0; 
    wire[6:0] frontend_tlb_must_alloc_array =7'h0; 
    wire[6:0] frontend_tlb_pf_st_array =7'h0; 
    wire[6:0] frontend_tlb_gf_ld_array =7'h0; 
    wire[6:0] frontend_tlb_gf_st_array =7'h0; 
    wire[6:0] frontend_tlb_gf_inst_array =7'h0; 
    wire[5:0] frontend_tlb_stage2_bypass =6'h3F; 
    wire[5:0] frontend_tlb_gpa_hits_hit_mask =6'h3F; 
    wire[5:0] frontend_tlb_gpa_hits =6'h3F; 
    wire[21:0] frontend_tlb_satp_ppn =22'h0; 
    wire[8:0] frontend_tlb_satp_asid =9'h0; 
    wire[19:0] frontend_tlb_vpn = frontend_tlb_io_req_bits_vaddr [31:12]; 
    wire[19:0] frontend_tlb_ppn = frontend_tlb_vpn ; 
    wire[19:0] frontend_tlb_refill_ppn = frontend_tlb_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire[19:0] frontend_tlb_newEntry_ppn = frontend_tlb_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire[19:0] frontend_tlb_mpu_ppn = frontend_tlb_io_req_bits_vaddr [31:12]; 
    wire[11:0] frontend_tlb_io_resp_gpa_offset = frontend_tlb_io_req_bits_vaddr [11:0]; 
    wire[31:0] frontend_tlb_mpu_physaddr ={ frontend_tlb_mpu_ppn , frontend_tlb_io_resp_gpa_offset }; 
    wire[2:0] frontend_tlb_mpu_priv ={ frontend_tlb_io_ptw_status_debug ,2'h3}; 
    wire[19:0] frontend_tlb__GEN ={ frontend_tlb_mpu_physaddr [31:14],~( frontend_tlb_mpu_physaddr [13:12])}; 
    wire[5:0] frontend_tlb__GEN_0 ={ frontend_tlb_mpu_physaddr [31:28],~( frontend_tlb_mpu_physaddr [27:26])}; 
    wire[9:0] frontend_tlb__GEN_1 = frontend_tlb_mpu_physaddr [25:16]^10'h200; 
    wire[15:0] frontend_tlb__GEN_2 ={ frontend_tlb_mpu_physaddr [31:26], frontend_tlb__GEN_1 }; 
    wire frontend_tlb__GEN_3 = frontend_tlb_mpu_physaddr [31:14]!=18'h20000; 
    wire[15:0] frontend_tlb__GEN_4 ={ frontend_tlb_mpu_physaddr [31:17],~( frontend_tlb_mpu_physaddr [16])}; 
    wire[2:0] frontend_tlb__GEN_5 ={ frontend_tlb_mpu_physaddr [31],~( frontend_tlb_mpu_physaddr [30:29])}; 
    wire frontend_tlb_legal_address =~(| frontend_tlb__GEN )|~(| frontend_tlb__GEN_0 )|~(| frontend_tlb__GEN_2 )|~ frontend_tlb__GEN_3 |~(|( frontend_tlb_mpu_physaddr [31:12]))|~(| frontend_tlb__GEN_4 )|~(| frontend_tlb__GEN_5 ); 
    wire frontend_tlb_homogeneous =~(|( frontend_tlb_mpu_physaddr [31:12]))|~(| frontend_tlb__GEN )|~(| frontend_tlb__GEN_4 )|~(| frontend_tlb__GEN_2 )|~(| frontend_tlb__GEN_0 )|~(| frontend_tlb__GEN_5 )|~ frontend_tlb__GEN_3 ; 
    wire frontend_tlb_deny_access_to_debug =~( frontend_tlb_mpu_priv [2])&~(|( frontend_tlb_mpu_physaddr [31:12])); 
    wire frontend_tlb_prot_r = frontend_tlb_legal_address &~ frontend_tlb_deny_access_to_debug & frontend_tlb__pmp_io_r ; 
    wire frontend_tlb_newEntry_pr = frontend_tlb_prot_r ; 
    wire[2:0] frontend_tlb__GEN_6 ={ frontend_tlb_mpu_physaddr [30], frontend_tlb_mpu_physaddr [27], frontend_tlb_mpu_physaddr [16]}; 
    wire[2:0] frontend_tlb__GEN_7 ={ frontend_tlb_mpu_physaddr [31:30],~( frontend_tlb_mpu_physaddr [27])}; 
    wire[1:0] frontend_tlb__GEN_8 ={ frontend_tlb_mpu_physaddr [31],~( frontend_tlb_mpu_physaddr [30])}; 
    wire frontend_tlb_prot_w = frontend_tlb_legal_address &(~(| frontend_tlb__GEN_6 )|~(| frontend_tlb__GEN_7 )|~(| frontend_tlb__GEN_8 ))&~ frontend_tlb_deny_access_to_debug & frontend_tlb__pmp_io_w ; 
    wire frontend_tlb_newEntry_pw = frontend_tlb_prot_w ; 
    wire frontend_tlb_prot_pp = frontend_tlb_legal_address &(~(| frontend_tlb__GEN_6 )|~(| frontend_tlb__GEN_7 )|~(| frontend_tlb__GEN_8 )); 
    wire frontend_tlb_newEntry_ppp = frontend_tlb_prot_pp ; 
    wire frontend_tlb_prot_al = frontend_tlb_legal_address &(~(| frontend_tlb__GEN_6 )|~(| frontend_tlb__GEN_7 )); 
    wire frontend_tlb_newEntry_pal = frontend_tlb_prot_al ; 
    wire frontend_tlb_prot_aa = frontend_tlb_legal_address &(~(| frontend_tlb__GEN_6 )|~(| frontend_tlb__GEN_7 )); 
    wire frontend_tlb_newEntry_paa = frontend_tlb_prot_aa ; 
    wire frontend_tlb_prot_x = frontend_tlb_legal_address &({ frontend_tlb_mpu_physaddr [30], frontend_tlb_mpu_physaddr [27], frontend_tlb_mpu_physaddr [25]}==3'h0|~(| frontend_tlb__GEN_8 ))&~ frontend_tlb_deny_access_to_debug & frontend_tlb__pmp_io_x ; 
    wire frontend_tlb_newEntry_px = frontend_tlb_prot_x ; 
    wire frontend_tlb_prot_eff = frontend_tlb_legal_address &({ frontend_tlb_mpu_physaddr [31:30], frontend_tlb_mpu_physaddr [27], frontend_tlb_mpu_physaddr [25], frontend_tlb_mpu_physaddr [16], frontend_tlb_mpu_physaddr [13]}==6'h0|{ frontend_tlb_mpu_physaddr [31:30], frontend_tlb_mpu_physaddr [27], frontend_tlb__GEN_1 [9], frontend_tlb_mpu_physaddr [16]}==5'h0|~(| frontend_tlb__GEN_7 )|~(| frontend_tlb__GEN_8 )); 
    wire frontend_tlb_newEntry_eff = frontend_tlb_prot_eff ; 
    wire[1:0] frontend_tlb_hitsVec_idx = frontend_tlb_vpn [1:0]; 
    wire frontend_tlb_newEntry_g = frontend_tlb_io_ptw_resp_bits_pte_g & frontend_tlb_io_ptw_resp_bits_pte_v ; 
    wire frontend_tlb_newEntry_sr = frontend_tlb_io_ptw_resp_bits_pte_v &( frontend_tlb_io_ptw_resp_bits_pte_r | frontend_tlb_io_ptw_resp_bits_pte_x &~ frontend_tlb_io_ptw_resp_bits_pte_w )& frontend_tlb_io_ptw_resp_bits_pte_a & frontend_tlb_io_ptw_resp_bits_pte_r ; 
    wire frontend_tlb_newEntry_sw = frontend_tlb_io_ptw_resp_bits_pte_v &( frontend_tlb_io_ptw_resp_bits_pte_r | frontend_tlb_io_ptw_resp_bits_pte_x &~ frontend_tlb_io_ptw_resp_bits_pte_w )& frontend_tlb_io_ptw_resp_bits_pte_a & frontend_tlb_io_ptw_resp_bits_pte_w & frontend_tlb_io_ptw_resp_bits_pte_d ; 
    wire frontend_tlb_newEntry_sx = frontend_tlb_io_ptw_resp_bits_pte_v &( frontend_tlb_io_ptw_resp_bits_pte_r | frontend_tlb_io_ptw_resp_bits_pte_x &~ frontend_tlb_io_ptw_resp_bits_pte_w )& frontend_tlb_io_ptw_resp_bits_pte_a & frontend_tlb_io_ptw_resp_bits_pte_x ; 
    wire[1:0] frontend_tlb__GEN_9 ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_lo_hi_hi ; 
  assign  frontend_tlb_special_entry_data_0_lo_lo_hi_hi = frontend_tlb__GEN_9 ; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_lo_lo_hi_hi = frontend_tlb__GEN_9 ; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_lo_lo_hi_hi = frontend_tlb__GEN_9 ; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_lo_lo_hi_hi = frontend_tlb__GEN_9 ; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_lo_lo_hi_hi = frontend_tlb__GEN_9 ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_lo_hi_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_lo_lo_hi_hi = frontend_tlb__GEN_9 ; 
    wire[2:0] frontend_tlb_special_entry_data_0_lo_lo_hi ={ frontend_tlb_special_entry_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_special_entry_data_0_lo_lo ={ frontend_tlb_special_entry_data_0_lo_lo_hi ,2'h0}; 
    wire[1:0] frontend_tlb__GEN_10 ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_hi_lo_hi ; 
  assign  frontend_tlb_special_entry_data_0_lo_hi_lo_hi = frontend_tlb__GEN_10 ; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_lo_hi_lo_hi = frontend_tlb__GEN_10 ; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_lo_hi_lo_hi = frontend_tlb__GEN_10 ; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_lo_hi_lo_hi = frontend_tlb__GEN_10 ; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_lo_hi_lo_hi = frontend_tlb__GEN_10 ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_lo_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_lo_hi_lo_hi = frontend_tlb__GEN_10 ; 
    wire[2:0] frontend_tlb_special_entry_data_0_lo_hi_lo ={ frontend_tlb_special_entry_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb__GEN_11 ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_hi_hi_hi ; 
  assign  frontend_tlb_special_entry_data_0_lo_hi_hi_hi = frontend_tlb__GEN_11 ; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_lo_hi_hi_hi = frontend_tlb__GEN_11 ; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_lo_hi_hi_hi = frontend_tlb__GEN_11 ; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_lo_hi_hi_hi = frontend_tlb__GEN_11 ; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_lo_hi_hi_hi = frontend_tlb__GEN_11 ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_hi_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_lo_hi_hi_hi = frontend_tlb__GEN_11 ; 
    wire[2:0] frontend_tlb_special_entry_data_0_lo_hi_hi ={ frontend_tlb_special_entry_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_special_entry_data_0_lo_hi ={ frontend_tlb_special_entry_data_0_lo_hi_hi , frontend_tlb_special_entry_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_special_entry_data_0_lo ={ frontend_tlb_special_entry_data_0_lo_hi , frontend_tlb_special_entry_data_0_lo_lo }; 
    wire[1:0] frontend_tlb__GEN_12 ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[1:0] frontend_tlb_special_entry_data_0_hi_lo_lo_hi ; 
  assign  frontend_tlb_special_entry_data_0_hi_lo_lo_hi = frontend_tlb__GEN_12 ; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_lo_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_hi_lo_lo_hi = frontend_tlb__GEN_12 ; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_lo_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_hi_lo_lo_hi = frontend_tlb__GEN_12 ; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_lo_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_hi_lo_lo_hi = frontend_tlb__GEN_12 ; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_lo_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_hi_lo_lo_hi = frontend_tlb__GEN_12 ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_lo_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_hi_lo_lo_hi = frontend_tlb__GEN_12 ; 
    wire[2:0] frontend_tlb_special_entry_data_0_hi_lo_lo ={ frontend_tlb_special_entry_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb__GEN_13 ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[1:0] frontend_tlb_special_entry_data_0_hi_lo_hi_hi ; 
  assign  frontend_tlb_special_entry_data_0_hi_lo_hi_hi = frontend_tlb__GEN_13 ; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_hi_lo_hi_hi = frontend_tlb__GEN_13 ; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_hi_lo_hi_hi = frontend_tlb__GEN_13 ; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_hi_lo_hi_hi = frontend_tlb__GEN_13 ; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_hi_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_hi_lo_hi_hi = frontend_tlb__GEN_13 ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_hi_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_hi_lo_hi_hi = frontend_tlb__GEN_13 ; 
    wire[2:0] frontend_tlb_special_entry_data_0_hi_lo_hi ={ frontend_tlb_special_entry_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_special_entry_data_0_hi_lo ={ frontend_tlb_special_entry_data_0_hi_lo_hi , frontend_tlb_special_entry_data_0_hi_lo_lo }; 
    wire[1:0] frontend_tlb__GEN_14 ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[1:0] frontend_tlb_special_entry_data_0_hi_hi_lo_hi ; 
  assign  frontend_tlb_special_entry_data_0_hi_hi_lo_hi = frontend_tlb__GEN_14 ; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_hi_hi_lo_hi = frontend_tlb__GEN_14 ; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_hi_hi_lo_hi = frontend_tlb__GEN_14 ; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_hi_hi_lo_hi = frontend_tlb__GEN_14 ; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_lo_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_hi_hi_lo_hi = frontend_tlb__GEN_14 ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_lo_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_hi_hi_lo_hi = frontend_tlb__GEN_14 ; 
    wire[2:0] frontend_tlb_special_entry_data_0_hi_hi_lo ={ frontend_tlb_special_entry_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb__GEN_15 ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[20:0] frontend_tlb_special_entry_data_0_hi_hi_hi_hi ; 
  assign  frontend_tlb_special_entry_data_0_hi_hi_hi_hi = frontend_tlb__GEN_15 ; 
    wire[20:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_0_data_0_hi_hi_hi_hi = frontend_tlb__GEN_15 ; 
    wire[20:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_1_data_0_hi_hi_hi_hi = frontend_tlb__GEN_15 ; 
    wire[20:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_2_data_0_hi_hi_hi_hi = frontend_tlb__GEN_15 ; 
    wire[20:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_hi_hi ; 
  assign  frontend_tlb_superpage_entries_3_data_0_hi_hi_hi_hi = frontend_tlb__GEN_15 ; 
    wire[20:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_hi_hi ; 
  assign  frontend_tlb_sectored_entries_0_0_data_hi_hi_hi_hi = frontend_tlb__GEN_15 ; 
    wire[21:0] frontend_tlb_special_entry_data_0_hi_hi_hi ={ frontend_tlb_special_entry_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_special_entry_data_0_hi_hi ={ frontend_tlb_special_entry_data_0_hi_hi_hi , frontend_tlb_special_entry_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_special_entry_data_0_hi ={ frontend_tlb_special_entry_data_0_hi_hi , frontend_tlb_special_entry_data_0_hi_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_0_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_0_data_0_lo_lo ={ frontend_tlb_superpage_entries_0_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_0_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_0_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_0_data_0_lo_hi ={ frontend_tlb_superpage_entries_0_data_0_lo_hi_hi , frontend_tlb_superpage_entries_0_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_0_data_0_lo ={ frontend_tlb_superpage_entries_0_data_0_lo_hi , frontend_tlb_superpage_entries_0_data_0_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_0_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_0_data_0_hi_lo ={ frontend_tlb_superpage_entries_0_data_0_hi_lo_hi , frontend_tlb_superpage_entries_0_data_0_hi_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_0_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[21:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_0_data_0_hi_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_hi_hi , frontend_tlb_superpage_entries_0_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_0_data_0_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_hi , frontend_tlb_superpage_entries_0_data_0_hi_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_1_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_1_data_0_lo_lo ={ frontend_tlb_superpage_entries_1_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_1_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_1_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_1_data_0_lo_hi ={ frontend_tlb_superpage_entries_1_data_0_lo_hi_hi , frontend_tlb_superpage_entries_1_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_1_data_0_lo ={ frontend_tlb_superpage_entries_1_data_0_lo_hi , frontend_tlb_superpage_entries_1_data_0_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_1_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_1_data_0_hi_lo ={ frontend_tlb_superpage_entries_1_data_0_hi_lo_hi , frontend_tlb_superpage_entries_1_data_0_hi_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_1_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[21:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_1_data_0_hi_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_hi_hi , frontend_tlb_superpage_entries_1_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_1_data_0_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_hi , frontend_tlb_superpage_entries_1_data_0_hi_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_2_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_2_data_0_lo_lo ={ frontend_tlb_superpage_entries_2_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_2_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_2_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_2_data_0_lo_hi ={ frontend_tlb_superpage_entries_2_data_0_lo_hi_hi , frontend_tlb_superpage_entries_2_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_2_data_0_lo ={ frontend_tlb_superpage_entries_2_data_0_lo_hi , frontend_tlb_superpage_entries_2_data_0_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_2_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_2_data_0_hi_lo ={ frontend_tlb_superpage_entries_2_data_0_hi_lo_hi , frontend_tlb_superpage_entries_2_data_0_hi_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_2_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[21:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_2_data_0_hi_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_hi_hi , frontend_tlb_superpage_entries_2_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_2_data_0_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_hi , frontend_tlb_superpage_entries_2_data_0_hi_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_3_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_3_data_0_lo_lo ={ frontend_tlb_superpage_entries_3_data_0_lo_lo_hi ,2'h0}; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_3_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_3_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_3_data_0_lo_hi ={ frontend_tlb_superpage_entries_3_data_0_lo_hi_hi , frontend_tlb_superpage_entries_3_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_3_data_0_lo ={ frontend_tlb_superpage_entries_3_data_0_lo_hi , frontend_tlb_superpage_entries_3_data_0_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_3_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_3_data_0_hi_lo ={ frontend_tlb_superpage_entries_3_data_0_hi_lo_hi , frontend_tlb_superpage_entries_3_data_0_hi_lo_lo }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_3_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[21:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_3_data_0_hi_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_hi_hi , frontend_tlb_superpage_entries_3_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_3_data_0_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_hi , frontend_tlb_superpage_entries_3_data_0_hi_lo }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_lo_lo_hi ={ frontend_tlb_sectored_entries_0_0_data_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_sectored_entries_0_0_data_lo_lo ={ frontend_tlb_sectored_entries_0_0_data_lo_lo_hi ,2'h0}; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_lo ={ frontend_tlb_sectored_entries_0_0_data_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_hi ={ frontend_tlb_sectored_entries_0_0_data_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_sectored_entries_0_0_data_lo_hi ={ frontend_tlb_sectored_entries_0_0_data_lo_hi_hi , frontend_tlb_sectored_entries_0_0_data_lo_hi_lo }; 
    wire[10:0] frontend_tlb_sectored_entries_0_0_data_lo ={ frontend_tlb_sectored_entries_0_0_data_lo_hi , frontend_tlb_sectored_entries_0_0_data_lo_lo }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_lo ={ frontend_tlb_sectored_entries_0_0_data_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_sectored_entries_0_0_data_hi_lo ={ frontend_tlb_sectored_entries_0_0_data_hi_lo_hi , frontend_tlb_sectored_entries_0_0_data_hi_lo_lo }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_lo ={ frontend_tlb_sectored_entries_0_0_data_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[21:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_sectored_entries_0_0_data_hi_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_hi_hi , frontend_tlb_sectored_entries_0_0_data_hi_hi_lo }; 
    wire[30:0] frontend_tlb_sectored_entries_0_0_data_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_hi , frontend_tlb_sectored_entries_0_0_data_hi_lo }; 
    wire[1:0] frontend_tlb_ptw_ae_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_ae_ptw , frontend_tlb__entries_barrier_1_io_y_ae_ptw }; 
    wire[2:0] frontend_tlb_ptw_ae_array_lo ={ frontend_tlb_ptw_ae_array_lo_hi , frontend_tlb__entries_barrier_io_y_ae_ptw }; 
    wire[1:0] frontend_tlb_ptw_ae_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_ae_ptw , frontend_tlb__entries_barrier_4_io_y_ae_ptw }; 
    wire[2:0] frontend_tlb_ptw_ae_array_hi ={ frontend_tlb_ptw_ae_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_ae_ptw }; 
    wire[6:0] frontend_tlb_ptw_ae_array ={1'h0, frontend_tlb_ptw_ae_array_hi , frontend_tlb_ptw_ae_array_lo }; 
    wire[1:0] frontend_tlb_final_ae_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_ae_final , frontend_tlb__entries_barrier_1_io_y_ae_final }; 
    wire[2:0] frontend_tlb_final_ae_array_lo ={ frontend_tlb_final_ae_array_lo_hi , frontend_tlb__entries_barrier_io_y_ae_final }; 
    wire[1:0] frontend_tlb_final_ae_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_ae_final , frontend_tlb__entries_barrier_4_io_y_ae_final }; 
    wire[2:0] frontend_tlb_final_ae_array_hi ={ frontend_tlb_final_ae_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_ae_final }; 
    wire[6:0] frontend_tlb_final_ae_array ={1'h0, frontend_tlb_final_ae_array_hi , frontend_tlb_final_ae_array_lo }; 
    wire[1:0] frontend_tlb_ptw_pf_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_pf , frontend_tlb__entries_barrier_1_io_y_pf }; 
    wire[2:0] frontend_tlb_ptw_pf_array_lo ={ frontend_tlb_ptw_pf_array_lo_hi , frontend_tlb__entries_barrier_io_y_pf }; 
    wire[1:0] frontend_tlb_ptw_pf_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_pf , frontend_tlb__entries_barrier_4_io_y_pf }; 
    wire[2:0] frontend_tlb_ptw_pf_array_hi ={ frontend_tlb_ptw_pf_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_pf }; 
    wire[6:0] frontend_tlb_ptw_pf_array ={1'h0, frontend_tlb_ptw_pf_array_hi , frontend_tlb_ptw_pf_array_lo }; 
    wire[1:0] frontend_tlb_ptw_gf_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_gf , frontend_tlb__entries_barrier_1_io_y_gf }; 
    wire[2:0] frontend_tlb_ptw_gf_array_lo ={ frontend_tlb_ptw_gf_array_lo_hi , frontend_tlb__entries_barrier_io_y_gf }; 
    wire[1:0] frontend_tlb_ptw_gf_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_gf , frontend_tlb__entries_barrier_4_io_y_gf }; 
    wire[2:0] frontend_tlb_ptw_gf_array_hi ={ frontend_tlb_ptw_gf_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_gf }; 
    wire[6:0] frontend_tlb_ptw_gf_array ={1'h0, frontend_tlb_ptw_gf_array_hi , frontend_tlb_ptw_gf_array_lo }; 
    wire[1:0] frontend_tlb__GEN_16 ={ frontend_tlb__entries_barrier_2_io_y_u , frontend_tlb__entries_barrier_1_io_y_u }; 
    wire[1:0] frontend_tlb_priv_rw_ok_lo_hi ; 
  assign  frontend_tlb_priv_rw_ok_lo_hi = frontend_tlb__GEN_16 ; 
    wire[1:0] frontend_tlb_priv_rw_ok_lo_hi_1 ; 
  assign  frontend_tlb_priv_rw_ok_lo_hi_1 = frontend_tlb__GEN_16 ; 
    wire[1:0] frontend_tlb_priv_x_ok_lo_hi ; 
  assign  frontend_tlb_priv_x_ok_lo_hi = frontend_tlb__GEN_16 ; 
    wire[1:0] frontend_tlb_priv_x_ok_lo_hi_1 ; 
  assign  frontend_tlb_priv_x_ok_lo_hi_1 = frontend_tlb__GEN_16 ; 
    wire[2:0] frontend_tlb_priv_rw_ok_lo ={ frontend_tlb_priv_rw_ok_lo_hi , frontend_tlb__entries_barrier_io_y_u }; 
    wire[1:0] frontend_tlb__GEN_17 ={ frontend_tlb__entries_barrier_5_io_y_u , frontend_tlb__entries_barrier_4_io_y_u }; 
    wire[1:0] frontend_tlb_priv_rw_ok_hi_hi ; 
  assign  frontend_tlb_priv_rw_ok_hi_hi = frontend_tlb__GEN_17 ; 
    wire[1:0] frontend_tlb_priv_rw_ok_hi_hi_1 ; 
  assign  frontend_tlb_priv_rw_ok_hi_hi_1 = frontend_tlb__GEN_17 ; 
    wire[1:0] frontend_tlb_priv_x_ok_hi_hi ; 
  assign  frontend_tlb_priv_x_ok_hi_hi = frontend_tlb__GEN_17 ; 
    wire[1:0] frontend_tlb_priv_x_ok_hi_hi_1 ; 
  assign  frontend_tlb_priv_x_ok_hi_hi_1 = frontend_tlb__GEN_17 ; 
    wire[2:0] frontend_tlb_priv_rw_ok_hi ={ frontend_tlb_priv_rw_ok_hi_hi , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[2:0] frontend_tlb_priv_rw_ok_lo_1 ={ frontend_tlb_priv_rw_ok_lo_hi_1 , frontend_tlb__entries_barrier_io_y_u }; 
    wire[2:0] frontend_tlb_priv_rw_ok_hi_1 ={ frontend_tlb_priv_rw_ok_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[5:0] frontend_tlb_priv_rw_ok =~{ frontend_tlb_priv_rw_ok_hi_1 , frontend_tlb_priv_rw_ok_lo_1 }; 
    wire[2:0] frontend_tlb_priv_x_ok_lo ={ frontend_tlb_priv_x_ok_lo_hi , frontend_tlb__entries_barrier_io_y_u }; 
    wire[2:0] frontend_tlb_priv_x_ok_hi ={ frontend_tlb_priv_x_ok_hi_hi , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[5:0] frontend_tlb_priv_x_ok =~{ frontend_tlb_priv_x_ok_hi , frontend_tlb_priv_x_ok_lo }; 
    wire[2:0] frontend_tlb_priv_x_ok_lo_1 ={ frontend_tlb_priv_x_ok_lo_hi_1 , frontend_tlb__entries_barrier_io_y_u }; 
    wire[2:0] frontend_tlb_priv_x_ok_hi_1 ={ frontend_tlb_priv_x_ok_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[1:0] frontend_tlb_stage1_bypass_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_ae_stage2 , frontend_tlb__entries_barrier_1_io_y_ae_stage2 }; 
    wire[2:0] frontend_tlb_stage1_bypass_lo ={ frontend_tlb_stage1_bypass_lo_hi , frontend_tlb__entries_barrier_io_y_ae_stage2 }; 
    wire[1:0] frontend_tlb_stage1_bypass_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_ae_stage2 , frontend_tlb__entries_barrier_4_io_y_ae_stage2 }; 
    wire[2:0] frontend_tlb_stage1_bypass_hi ={ frontend_tlb_stage1_bypass_hi_hi , frontend_tlb__entries_barrier_3_io_y_ae_stage2 }; 
    wire[1:0] frontend_tlb_r_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_sr , frontend_tlb__entries_barrier_1_io_y_sr }; 
    wire[2:0] frontend_tlb_r_array_lo ={ frontend_tlb_r_array_lo_hi , frontend_tlb__entries_barrier_io_y_sr }; 
    wire[1:0] frontend_tlb_r_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_sr , frontend_tlb__entries_barrier_4_io_y_sr }; 
    wire[2:0] frontend_tlb_r_array_hi ={ frontend_tlb_r_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_sr }; 
    wire[1:0] frontend_tlb__GEN_18 ={ frontend_tlb__entries_barrier_2_io_y_sx , frontend_tlb__entries_barrier_1_io_y_sx }; 
    wire[1:0] frontend_tlb_r_array_lo_hi_1 ; 
  assign  frontend_tlb_r_array_lo_hi_1 = frontend_tlb__GEN_18 ; 
    wire[1:0] frontend_tlb_x_array_lo_hi ; 
  assign  frontend_tlb_x_array_lo_hi = frontend_tlb__GEN_18 ; 
    wire[2:0] frontend_tlb_r_array_lo_1 ={ frontend_tlb_r_array_lo_hi_1 , frontend_tlb__entries_barrier_io_y_sx }; 
    wire[1:0] frontend_tlb__GEN_19 ={ frontend_tlb__entries_barrier_5_io_y_sx , frontend_tlb__entries_barrier_4_io_y_sx }; 
    wire[1:0] frontend_tlb_r_array_hi_hi_1 ; 
  assign  frontend_tlb_r_array_hi_hi_1 = frontend_tlb__GEN_19 ; 
    wire[1:0] frontend_tlb_x_array_hi_hi ; 
  assign  frontend_tlb_x_array_hi_hi = frontend_tlb__GEN_19 ; 
    wire[2:0] frontend_tlb_r_array_hi_1 ={ frontend_tlb_r_array_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_sx }; 
    wire[6:0] frontend_tlb_r_array ={1'h1, frontend_tlb_priv_rw_ok &{ frontend_tlb_r_array_hi , frontend_tlb_r_array_lo }}; 
    wire[1:0] frontend_tlb_w_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_sw , frontend_tlb__entries_barrier_1_io_y_sw }; 
    wire[2:0] frontend_tlb_w_array_lo ={ frontend_tlb_w_array_lo_hi , frontend_tlb__entries_barrier_io_y_sw }; 
    wire[1:0] frontend_tlb_w_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_sw , frontend_tlb__entries_barrier_4_io_y_sw }; 
    wire[2:0] frontend_tlb_w_array_hi ={ frontend_tlb_w_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_sw }; 
    wire[6:0] frontend_tlb_w_array ={1'h1, frontend_tlb_priv_rw_ok &{ frontend_tlb_w_array_hi , frontend_tlb_w_array_lo }}; 
    wire[2:0] frontend_tlb_x_array_lo ={ frontend_tlb_x_array_lo_hi , frontend_tlb__entries_barrier_io_y_sx }; 
    wire[2:0] frontend_tlb_x_array_hi ={ frontend_tlb_x_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_sx }; 
    wire[6:0] frontend_tlb_x_array ={1'h1, frontend_tlb_priv_x_ok &{ frontend_tlb_x_array_hi , frontend_tlb_x_array_lo }}; 
    wire[1:0] frontend_tlb_hr_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_hr , frontend_tlb__entries_barrier_1_io_y_hr }; 
    wire[2:0] frontend_tlb_hr_array_lo ={ frontend_tlb_hr_array_lo_hi , frontend_tlb__entries_barrier_io_y_hr }; 
    wire[1:0] frontend_tlb_hr_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_hr , frontend_tlb__entries_barrier_4_io_y_hr }; 
    wire[2:0] frontend_tlb_hr_array_hi ={ frontend_tlb_hr_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_hr }; 
    wire[1:0] frontend_tlb__GEN_20 ={ frontend_tlb__entries_barrier_2_io_y_hx , frontend_tlb__entries_barrier_1_io_y_hx }; 
    wire[1:0] frontend_tlb_hr_array_lo_hi_1 ; 
  assign  frontend_tlb_hr_array_lo_hi_1 = frontend_tlb__GEN_20 ; 
    wire[1:0] frontend_tlb_hx_array_lo_hi ; 
  assign  frontend_tlb_hx_array_lo_hi = frontend_tlb__GEN_20 ; 
    wire[2:0] frontend_tlb_hr_array_lo_1 ={ frontend_tlb_hr_array_lo_hi_1 , frontend_tlb__entries_barrier_io_y_hx }; 
    wire[1:0] frontend_tlb__GEN_21 ={ frontend_tlb__entries_barrier_5_io_y_hx , frontend_tlb__entries_barrier_4_io_y_hx }; 
    wire[1:0] frontend_tlb_hr_array_hi_hi_1 ; 
  assign  frontend_tlb_hr_array_hi_hi_1 = frontend_tlb__GEN_21 ; 
    wire[1:0] frontend_tlb_hx_array_hi_hi ; 
  assign  frontend_tlb_hx_array_hi_hi = frontend_tlb__GEN_21 ; 
    wire[2:0] frontend_tlb_hr_array_hi_1 ={ frontend_tlb_hr_array_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_hx }; 
    wire[1:0] frontend_tlb_hw_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_hw , frontend_tlb__entries_barrier_1_io_y_hw }; 
    wire[2:0] frontend_tlb_hw_array_lo ={ frontend_tlb_hw_array_lo_hi , frontend_tlb__entries_barrier_io_y_hw }; 
    wire[1:0] frontend_tlb_hw_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_hw , frontend_tlb__entries_barrier_4_io_y_hw }; 
    wire[2:0] frontend_tlb_hw_array_hi ={ frontend_tlb_hw_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_hw }; 
    wire[2:0] frontend_tlb_hx_array_lo ={ frontend_tlb_hx_array_lo_hi , frontend_tlb__entries_barrier_io_y_hx }; 
    wire[2:0] frontend_tlb_hx_array_hi ={ frontend_tlb_hx_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_hx }; 
    wire[1:0] frontend_tlb_pr_array_lo ={ frontend_tlb__entries_barrier_1_io_y_pr , frontend_tlb__entries_barrier_io_y_pr }; 
    wire[1:0] frontend_tlb_pr_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_pr , frontend_tlb__entries_barrier_3_io_y_pr }; 
    wire[2:0] frontend_tlb_pr_array_hi ={ frontend_tlb_pr_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_pr }; 
    wire[6:0] frontend_tlb__px_array_T_4 = frontend_tlb_ptw_ae_array | frontend_tlb_final_ae_array ; 
    wire[6:0] frontend_tlb_pr_array ={{2{ frontend_tlb_prot_r }}, frontend_tlb_pr_array_hi , frontend_tlb_pr_array_lo }&~ frontend_tlb__px_array_T_4 ; 
    wire[1:0] frontend_tlb_pw_array_lo ={ frontend_tlb__entries_barrier_1_io_y_pw , frontend_tlb__entries_barrier_io_y_pw }; 
    wire[1:0] frontend_tlb_pw_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_pw , frontend_tlb__entries_barrier_3_io_y_pw }; 
    wire[2:0] frontend_tlb_pw_array_hi ={ frontend_tlb_pw_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_pw }; 
    wire[6:0] frontend_tlb_pw_array ={{2{ frontend_tlb_prot_w }}, frontend_tlb_pw_array_hi , frontend_tlb_pw_array_lo }&~ frontend_tlb__px_array_T_4 ; 
    wire[1:0] frontend_tlb_px_array_lo ={ frontend_tlb__entries_barrier_1_io_y_px , frontend_tlb__entries_barrier_io_y_px }; 
    wire[1:0] frontend_tlb_px_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_px , frontend_tlb__entries_barrier_3_io_y_px }; 
    wire[2:0] frontend_tlb_px_array_hi ={ frontend_tlb_px_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_px }; 
    wire[6:0] frontend_tlb_px_array ={{2{ frontend_tlb_prot_x }}, frontend_tlb_px_array_hi , frontend_tlb_px_array_lo }&~ frontend_tlb__px_array_T_4 ; 
    wire[1:0] frontend_tlb_eff_array_lo ={ frontend_tlb__entries_barrier_1_io_y_eff , frontend_tlb__entries_barrier_io_y_eff }; 
    wire[1:0] frontend_tlb_eff_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_eff , frontend_tlb__entries_barrier_3_io_y_eff }; 
    wire[2:0] frontend_tlb_eff_array_hi ={ frontend_tlb_eff_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_eff }; 
    wire[6:0] frontend_tlb_eff_array ={{2{ frontend_tlb_prot_eff }}, frontend_tlb_eff_array_hi , frontend_tlb_eff_array_lo }; 
    wire[1:0] frontend_tlb__GEN_22 ={ frontend_tlb__entries_barrier_1_io_y_c , frontend_tlb__entries_barrier_io_y_c }; 
    wire[1:0] frontend_tlb_c_array_lo ; 
  assign  frontend_tlb_c_array_lo = frontend_tlb__GEN_22 ; 
    wire[1:0] frontend_tlb_prefetchable_array_lo ; 
  assign  frontend_tlb_prefetchable_array_lo = frontend_tlb__GEN_22 ; 
    wire[1:0] frontend_tlb__GEN_23 ={ frontend_tlb__entries_barrier_4_io_y_c , frontend_tlb__entries_barrier_3_io_y_c }; 
    wire[1:0] frontend_tlb_c_array_hi_hi ; 
  assign  frontend_tlb_c_array_hi_hi = frontend_tlb__GEN_23 ; 
    wire[1:0] frontend_tlb_prefetchable_array_hi_hi ; 
  assign  frontend_tlb_prefetchable_array_hi_hi = frontend_tlb__GEN_23 ; 
    wire[2:0] frontend_tlb_c_array_hi ={ frontend_tlb_c_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_c }; 
    wire[6:0] frontend_tlb_c_array ={2'h0, frontend_tlb_c_array_hi , frontend_tlb_c_array_lo }; 
    wire[1:0] frontend_tlb_ppp_array_lo ={ frontend_tlb__entries_barrier_1_io_y_ppp , frontend_tlb__entries_barrier_io_y_ppp }; 
    wire[1:0] frontend_tlb_ppp_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_ppp , frontend_tlb__entries_barrier_3_io_y_ppp }; 
    wire[2:0] frontend_tlb_ppp_array_hi ={ frontend_tlb_ppp_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_ppp }; 
    wire[6:0] frontend_tlb_ppp_array ={{2{ frontend_tlb_prot_pp }}, frontend_tlb_ppp_array_hi , frontend_tlb_ppp_array_lo }; 
    wire[1:0] frontend_tlb_paa_array_lo ={ frontend_tlb__entries_barrier_1_io_y_paa , frontend_tlb__entries_barrier_io_y_paa }; 
    wire[1:0] frontend_tlb_paa_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_paa , frontend_tlb__entries_barrier_3_io_y_paa }; 
    wire[2:0] frontend_tlb_paa_array_hi ={ frontend_tlb_paa_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_paa }; 
    wire[6:0] frontend_tlb_paa_array ={{2{ frontend_tlb_prot_aa }}, frontend_tlb_paa_array_hi , frontend_tlb_paa_array_lo }; 
    wire[1:0] frontend_tlb_pal_array_lo ={ frontend_tlb__entries_barrier_1_io_y_pal , frontend_tlb__entries_barrier_io_y_pal }; 
    wire[1:0] frontend_tlb_pal_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_pal , frontend_tlb__entries_barrier_3_io_y_pal }; 
    wire[2:0] frontend_tlb_pal_array_hi ={ frontend_tlb_pal_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_pal }; 
    wire[6:0] frontend_tlb_pal_array ={{2{ frontend_tlb_prot_al }}, frontend_tlb_pal_array_hi , frontend_tlb_pal_array_lo }; 
    wire[6:0] frontend_tlb_ppp_array_if_cached = frontend_tlb_ppp_array | frontend_tlb_c_array ; 
    wire[6:0] frontend_tlb_paa_array_if_cached = frontend_tlb_paa_array | frontend_tlb_c_array ; 
    wire[6:0] frontend_tlb_pal_array_if_cached = frontend_tlb_pal_array | frontend_tlb_c_array ; 
    wire[2:0] frontend_tlb_prefetchable_array_hi ={ frontend_tlb_prefetchable_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_c }; 
    wire[6:0] frontend_tlb_prefetchable_array ={2'h0, frontend_tlb_prefetchable_array_hi , frontend_tlb_prefetchable_array_lo }; 
    wire frontend_tlb_misaligned =|( frontend_tlb_io_req_bits_vaddr [1:0]); 
    wire[6:0] frontend_tlb_ae_array = frontend_tlb_misaligned  ?  frontend_tlb_eff_array :7'h0; 
    wire[6:0] frontend_tlb_ae_ld_array = frontend_tlb_ae_array |~ frontend_tlb_pr_array ; 
    wire[6:0] frontend_tlb_pf_ld_array =(~ frontend_tlb_r_array &~ frontend_tlb_ptw_ae_array | frontend_tlb_ptw_pf_array )&~ frontend_tlb_ptw_gf_array ; 
    wire[6:0] frontend_tlb_pf_inst_array =(~ frontend_tlb_x_array &~ frontend_tlb_ptw_ae_array | frontend_tlb_ptw_pf_array )&~ frontend_tlb_ptw_gf_array ; 
    wire[1:0] frontend_tlb_lo ={ frontend_tlb_superpage_hits_1 , frontend_tlb_superpage_hits_0 }; 
    wire[1:0] frontend_tlb_lo_1 = frontend_tlb_lo ; 
    wire[1:0] frontend_tlb_hi ={ frontend_tlb_superpage_hits_3 , frontend_tlb_superpage_hits_2 }; 
    wire[1:0] frontend_tlb_hi_1 = frontend_tlb_hi ; 
    wire[1:0] frontend_tlb_state_reg_touch_way_sized ={| frontend_tlb_hi_1 , frontend_tlb_hi_1 [1]| frontend_tlb_lo_1 [1]}; 
    wire frontend_tlb_state_reg_set_left_older =~( frontend_tlb_state_reg_touch_way_sized [1]); 
    wire[1:0] frontend_tlb_state_reg_hi ={ frontend_tlb_state_reg_set_left_older ,~ frontend_tlb_state_reg_set_left_older &~( frontend_tlb_state_reg_touch_way_sized [0])}; 
    wire[20:0] frontend_tlb_io_resp_gpa_page ={1'h0, frontend_tlb_vpn };  
    wire[1:0] frontend_tlb_pmp_io_prv;
    wire frontend_tlb_pmp_io_pmp_0_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_0_cfg_a;
    wire frontend_tlb_pmp_io_pmp_0_cfg_x;
    wire frontend_tlb_pmp_io_pmp_0_cfg_w;
    wire frontend_tlb_pmp_io_pmp_0_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_0_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_0_mask;
    wire frontend_tlb_pmp_io_pmp_1_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_1_cfg_a;
    wire frontend_tlb_pmp_io_pmp_1_cfg_x;
    wire frontend_tlb_pmp_io_pmp_1_cfg_w;
    wire frontend_tlb_pmp_io_pmp_1_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_1_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_1_mask;
    wire frontend_tlb_pmp_io_pmp_2_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_2_cfg_a;
    wire frontend_tlb_pmp_io_pmp_2_cfg_x;
    wire frontend_tlb_pmp_io_pmp_2_cfg_w;
    wire frontend_tlb_pmp_io_pmp_2_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_2_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_2_mask;
    wire frontend_tlb_pmp_io_pmp_3_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_3_cfg_a;
    wire frontend_tlb_pmp_io_pmp_3_cfg_x;
    wire frontend_tlb_pmp_io_pmp_3_cfg_w;
    wire frontend_tlb_pmp_io_pmp_3_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_3_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_3_mask;
    wire frontend_tlb_pmp_io_pmp_4_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_4_cfg_a;
    wire frontend_tlb_pmp_io_pmp_4_cfg_x;
    wire frontend_tlb_pmp_io_pmp_4_cfg_w;
    wire frontend_tlb_pmp_io_pmp_4_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_4_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_4_mask;
    wire frontend_tlb_pmp_io_pmp_5_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_5_cfg_a;
    wire frontend_tlb_pmp_io_pmp_5_cfg_x;
    wire frontend_tlb_pmp_io_pmp_5_cfg_w;
    wire frontend_tlb_pmp_io_pmp_5_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_5_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_5_mask;
    wire frontend_tlb_pmp_io_pmp_6_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_6_cfg_a;
    wire frontend_tlb_pmp_io_pmp_6_cfg_x;
    wire frontend_tlb_pmp_io_pmp_6_cfg_w;
    wire frontend_tlb_pmp_io_pmp_6_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_6_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_6_mask;
    wire frontend_tlb_pmp_io_pmp_7_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_7_cfg_a;
    wire frontend_tlb_pmp_io_pmp_7_cfg_x;
    wire frontend_tlb_pmp_io_pmp_7_cfg_w;
    wire frontend_tlb_pmp_io_pmp_7_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_7_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_7_mask;
    wire[31:0] frontend_tlb_pmp_io_addr;
    wire frontend_tlb_pmp_io_r;
    wire frontend_tlb_pmp_io_w;
    wire frontend_tlb_pmp_io_x;

    wire frontend_tlb_pmp_res_cur_cfg_l = frontend_tlb_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_cfg_a = frontend_tlb_pmp_io_pmp_7_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_addr = frontend_tlb_pmp_io_pmp_7_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_mask = frontend_tlb_pmp_io_pmp_7_mask ; 
    wire frontend_tlb_pmp_res_cur_1_cfg_l = frontend_tlb_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_1_cfg_a = frontend_tlb_pmp_io_pmp_6_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_1_addr = frontend_tlb_pmp_io_pmp_6_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_1_mask = frontend_tlb_pmp_io_pmp_6_mask ; 
    wire frontend_tlb_pmp_res_cur_2_cfg_l = frontend_tlb_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_2_cfg_a = frontend_tlb_pmp_io_pmp_5_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_2_addr = frontend_tlb_pmp_io_pmp_5_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_2_mask = frontend_tlb_pmp_io_pmp_5_mask ; 
    wire frontend_tlb_pmp_res_cur_3_cfg_l = frontend_tlb_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_3_cfg_a = frontend_tlb_pmp_io_pmp_4_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_3_addr = frontend_tlb_pmp_io_pmp_4_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_3_mask = frontend_tlb_pmp_io_pmp_4_mask ; 
    wire frontend_tlb_pmp_res_cur_4_cfg_l = frontend_tlb_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_4_cfg_a = frontend_tlb_pmp_io_pmp_3_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_4_addr = frontend_tlb_pmp_io_pmp_3_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_4_mask = frontend_tlb_pmp_io_pmp_3_mask ; 
    wire frontend_tlb_pmp_res_cur_5_cfg_l = frontend_tlb_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_5_cfg_a = frontend_tlb_pmp_io_pmp_2_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_5_addr = frontend_tlb_pmp_io_pmp_2_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_5_mask = frontend_tlb_pmp_io_pmp_2_mask ; 
    wire frontend_tlb_pmp_res_cur_6_cfg_l = frontend_tlb_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_6_cfg_a = frontend_tlb_pmp_io_pmp_1_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_6_addr = frontend_tlb_pmp_io_pmp_1_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_6_mask = frontend_tlb_pmp_io_pmp_1_mask ; 
    wire frontend_tlb_pmp_res_cur_7_cfg_l = frontend_tlb_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_7_cfg_a = frontend_tlb_pmp_io_pmp_0_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_7_addr = frontend_tlb_pmp_io_pmp_0_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_7_mask = frontend_tlb_pmp_io_pmp_0_mask ; 
    wire[1:0] frontend_tlb_pmp_pmp0_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_pmp0_cfg_a =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_1_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_2_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_3_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_4_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_5_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_6_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cur_7_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp_res_cfg_res =2'h0; 
    wire frontend_tlb_pmp_pmp0_cfg_l =1'h0; 
    wire[29:0] frontend_tlb_pmp_pmp0_addr =30'h0; 
    wire[31:0] frontend_tlb_pmp_pmp0_mask =32'h0; 
    wire frontend_tlb_pmp_default_0 = frontend_tlb_pmp_io_prv [1]; 
    wire frontend_tlb_pmp_pmp0_cfg_x = frontend_tlb_pmp_default_0 ; 
    wire frontend_tlb_pmp_pmp0_cfg_w = frontend_tlb_pmp_default_0 ; 
    wire frontend_tlb_pmp_pmp0_cfg_r = frontend_tlb_pmp_default_0 ; 
    wire frontend_tlb_pmp_res_hit = frontend_tlb_pmp_io_pmp_7_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_7_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_7_mask )==32'h0: frontend_tlb_pmp_io_pmp_7_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_6_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_7_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi ; 
  assign  frontend_tlb_pmp_res_hi = frontend_tlb_pmp__GEN ; 
    wire[1:0] frontend_tlb_pmp_res_hi_1 ; 
  assign  frontend_tlb_pmp_res_hi_1 = frontend_tlb_pmp__GEN ; 
    wire[1:0] frontend_tlb_pmp_res_hi_2 ; 
  assign  frontend_tlb_pmp_res_hi_2 = frontend_tlb_pmp__GEN ; 
    wire[1:0] frontend_tlb_pmp_res_hi_3 ; 
  assign  frontend_tlb_pmp_res_hi_3 = frontend_tlb_pmp__GEN ; 
    wire[1:0] frontend_tlb_pmp_res_hi_4 ; 
  assign  frontend_tlb_pmp_res_hi_4 = frontend_tlb_pmp__GEN ; 
    wire[1:0] frontend_tlb_pmp_res_hi_5 ; 
  assign  frontend_tlb_pmp_res_hi_5 = frontend_tlb_pmp__GEN ; 
    wire frontend_tlb_pmp_res_cur_cfg_r = frontend_tlb_pmp_io_pmp_7_cfg_r | frontend_tlb_pmp_res_ignore ; 
    wire frontend_tlb_pmp_res_cur_cfg_w = frontend_tlb_pmp_io_pmp_7_cfg_w | frontend_tlb_pmp_res_ignore ; 
    wire frontend_tlb_pmp_res_cur_cfg_x = frontend_tlb_pmp_io_pmp_7_cfg_x | frontend_tlb_pmp_res_ignore ; 
    wire frontend_tlb_pmp_res_hit_1 = frontend_tlb_pmp_io_pmp_6_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_6_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_6_mask )==32'h0: frontend_tlb_pmp_io_pmp_6_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_5_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_6_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_1 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_0 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_6 ; 
  assign  frontend_tlb_pmp_res_hi_6 = frontend_tlb_pmp__GEN_0 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_7 ; 
  assign  frontend_tlb_pmp_res_hi_7 = frontend_tlb_pmp__GEN_0 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_8 ; 
  assign  frontend_tlb_pmp_res_hi_8 = frontend_tlb_pmp__GEN_0 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_9 ; 
  assign  frontend_tlb_pmp_res_hi_9 = frontend_tlb_pmp__GEN_0 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_10 ; 
  assign  frontend_tlb_pmp_res_hi_10 = frontend_tlb_pmp__GEN_0 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_11 ; 
  assign  frontend_tlb_pmp_res_hi_11 = frontend_tlb_pmp__GEN_0 ; 
    wire frontend_tlb_pmp_res_cur_1_cfg_r = frontend_tlb_pmp_io_pmp_6_cfg_r | frontend_tlb_pmp_res_ignore_1 ; 
    wire frontend_tlb_pmp_res_cur_1_cfg_w = frontend_tlb_pmp_io_pmp_6_cfg_w | frontend_tlb_pmp_res_ignore_1 ; 
    wire frontend_tlb_pmp_res_cur_1_cfg_x = frontend_tlb_pmp_io_pmp_6_cfg_x | frontend_tlb_pmp_res_ignore_1 ; 
    wire frontend_tlb_pmp_res_hit_2 = frontend_tlb_pmp_io_pmp_5_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_5_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_5_mask )==32'h0: frontend_tlb_pmp_io_pmp_5_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_4_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_5_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_2 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_1 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_12 ; 
  assign  frontend_tlb_pmp_res_hi_12 = frontend_tlb_pmp__GEN_1 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_13 ; 
  assign  frontend_tlb_pmp_res_hi_13 = frontend_tlb_pmp__GEN_1 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_14 ; 
  assign  frontend_tlb_pmp_res_hi_14 = frontend_tlb_pmp__GEN_1 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_15 ; 
  assign  frontend_tlb_pmp_res_hi_15 = frontend_tlb_pmp__GEN_1 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_16 ; 
  assign  frontend_tlb_pmp_res_hi_16 = frontend_tlb_pmp__GEN_1 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_17 ; 
  assign  frontend_tlb_pmp_res_hi_17 = frontend_tlb_pmp__GEN_1 ; 
    wire frontend_tlb_pmp_res_cur_2_cfg_r = frontend_tlb_pmp_io_pmp_5_cfg_r | frontend_tlb_pmp_res_ignore_2 ; 
    wire frontend_tlb_pmp_res_cur_2_cfg_w = frontend_tlb_pmp_io_pmp_5_cfg_w | frontend_tlb_pmp_res_ignore_2 ; 
    wire frontend_tlb_pmp_res_cur_2_cfg_x = frontend_tlb_pmp_io_pmp_5_cfg_x | frontend_tlb_pmp_res_ignore_2 ; 
    wire frontend_tlb_pmp_res_hit_3 = frontend_tlb_pmp_io_pmp_4_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_4_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_4_mask )==32'h0: frontend_tlb_pmp_io_pmp_4_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_3_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_4_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_3 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_2 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_18 ; 
  assign  frontend_tlb_pmp_res_hi_18 = frontend_tlb_pmp__GEN_2 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_19 ; 
  assign  frontend_tlb_pmp_res_hi_19 = frontend_tlb_pmp__GEN_2 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_20 ; 
  assign  frontend_tlb_pmp_res_hi_20 = frontend_tlb_pmp__GEN_2 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_21 ; 
  assign  frontend_tlb_pmp_res_hi_21 = frontend_tlb_pmp__GEN_2 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_22 ; 
  assign  frontend_tlb_pmp_res_hi_22 = frontend_tlb_pmp__GEN_2 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_23 ; 
  assign  frontend_tlb_pmp_res_hi_23 = frontend_tlb_pmp__GEN_2 ; 
    wire frontend_tlb_pmp_res_cur_3_cfg_r = frontend_tlb_pmp_io_pmp_4_cfg_r | frontend_tlb_pmp_res_ignore_3 ; 
    wire frontend_tlb_pmp_res_cur_3_cfg_w = frontend_tlb_pmp_io_pmp_4_cfg_w | frontend_tlb_pmp_res_ignore_3 ; 
    wire frontend_tlb_pmp_res_cur_3_cfg_x = frontend_tlb_pmp_io_pmp_4_cfg_x | frontend_tlb_pmp_res_ignore_3 ; 
    wire frontend_tlb_pmp_res_hit_4 = frontend_tlb_pmp_io_pmp_3_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_3_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_3_mask )==32'h0: frontend_tlb_pmp_io_pmp_3_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_2_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_3_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_4 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_3 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_24 ; 
  assign  frontend_tlb_pmp_res_hi_24 = frontend_tlb_pmp__GEN_3 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_25 ; 
  assign  frontend_tlb_pmp_res_hi_25 = frontend_tlb_pmp__GEN_3 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_26 ; 
  assign  frontend_tlb_pmp_res_hi_26 = frontend_tlb_pmp__GEN_3 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_27 ; 
  assign  frontend_tlb_pmp_res_hi_27 = frontend_tlb_pmp__GEN_3 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_28 ; 
  assign  frontend_tlb_pmp_res_hi_28 = frontend_tlb_pmp__GEN_3 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_29 ; 
  assign  frontend_tlb_pmp_res_hi_29 = frontend_tlb_pmp__GEN_3 ; 
    wire frontend_tlb_pmp_res_cur_4_cfg_r = frontend_tlb_pmp_io_pmp_3_cfg_r | frontend_tlb_pmp_res_ignore_4 ; 
    wire frontend_tlb_pmp_res_cur_4_cfg_w = frontend_tlb_pmp_io_pmp_3_cfg_w | frontend_tlb_pmp_res_ignore_4 ; 
    wire frontend_tlb_pmp_res_cur_4_cfg_x = frontend_tlb_pmp_io_pmp_3_cfg_x | frontend_tlb_pmp_res_ignore_4 ; 
    wire frontend_tlb_pmp_res_hit_5 = frontend_tlb_pmp_io_pmp_2_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_2_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_2_mask )==32'h0: frontend_tlb_pmp_io_pmp_2_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_1_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_2_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_5 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_4 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_30 ; 
  assign  frontend_tlb_pmp_res_hi_30 = frontend_tlb_pmp__GEN_4 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_31 ; 
  assign  frontend_tlb_pmp_res_hi_31 = frontend_tlb_pmp__GEN_4 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_32 ; 
  assign  frontend_tlb_pmp_res_hi_32 = frontend_tlb_pmp__GEN_4 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_33 ; 
  assign  frontend_tlb_pmp_res_hi_33 = frontend_tlb_pmp__GEN_4 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_34 ; 
  assign  frontend_tlb_pmp_res_hi_34 = frontend_tlb_pmp__GEN_4 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_35 ; 
  assign  frontend_tlb_pmp_res_hi_35 = frontend_tlb_pmp__GEN_4 ; 
    wire frontend_tlb_pmp_res_cur_5_cfg_r = frontend_tlb_pmp_io_pmp_2_cfg_r | frontend_tlb_pmp_res_ignore_5 ; 
    wire frontend_tlb_pmp_res_cur_5_cfg_w = frontend_tlb_pmp_io_pmp_2_cfg_w | frontend_tlb_pmp_res_ignore_5 ; 
    wire frontend_tlb_pmp_res_cur_5_cfg_x = frontend_tlb_pmp_io_pmp_2_cfg_x | frontend_tlb_pmp_res_ignore_5 ; 
    wire frontend_tlb_pmp_res_hit_6 = frontend_tlb_pmp_io_pmp_1_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_1_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_1_mask )==32'h0: frontend_tlb_pmp_io_pmp_1_cfg_a [0]& frontend_tlb_pmp_io_addr >={ frontend_tlb_pmp_io_pmp_0_addr ,2'h0}& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_1_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_6 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_5 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_36 ; 
  assign  frontend_tlb_pmp_res_hi_36 = frontend_tlb_pmp__GEN_5 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_37 ; 
  assign  frontend_tlb_pmp_res_hi_37 = frontend_tlb_pmp__GEN_5 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_38 ; 
  assign  frontend_tlb_pmp_res_hi_38 = frontend_tlb_pmp__GEN_5 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_39 ; 
  assign  frontend_tlb_pmp_res_hi_39 = frontend_tlb_pmp__GEN_5 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_40 ; 
  assign  frontend_tlb_pmp_res_hi_40 = frontend_tlb_pmp__GEN_5 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_41 ; 
  assign  frontend_tlb_pmp_res_hi_41 = frontend_tlb_pmp__GEN_5 ; 
    wire frontend_tlb_pmp_res_cur_6_cfg_r = frontend_tlb_pmp_io_pmp_1_cfg_r | frontend_tlb_pmp_res_ignore_6 ; 
    wire frontend_tlb_pmp_res_cur_6_cfg_w = frontend_tlb_pmp_io_pmp_1_cfg_w | frontend_tlb_pmp_res_ignore_6 ; 
    wire frontend_tlb_pmp_res_cur_6_cfg_x = frontend_tlb_pmp_io_pmp_1_cfg_x | frontend_tlb_pmp_res_ignore_6 ; 
    wire frontend_tlb_pmp_res_hit_7 = frontend_tlb_pmp_io_pmp_0_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^{ frontend_tlb_pmp_io_pmp_0_addr ,2'h0})&~ frontend_tlb_pmp_io_pmp_0_mask )==32'h0: frontend_tlb_pmp_io_pmp_0_cfg_a [0]& frontend_tlb_pmp_io_addr <{ frontend_tlb_pmp_io_pmp_0_addr ,2'h0}; 
    wire frontend_tlb_pmp_res_ignore_7 = frontend_tlb_pmp_default_0 &~ frontend_tlb_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] frontend_tlb_pmp__GEN_6 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_42 ; 
  assign  frontend_tlb_pmp_res_hi_42 = frontend_tlb_pmp__GEN_6 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_43 ; 
  assign  frontend_tlb_pmp_res_hi_43 = frontend_tlb_pmp__GEN_6 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_44 ; 
  assign  frontend_tlb_pmp_res_hi_44 = frontend_tlb_pmp__GEN_6 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_45 ; 
  assign  frontend_tlb_pmp_res_hi_45 = frontend_tlb_pmp__GEN_6 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_46 ; 
  assign  frontend_tlb_pmp_res_hi_46 = frontend_tlb_pmp__GEN_6 ; 
    wire[1:0] frontend_tlb_pmp_res_hi_47 ; 
  assign  frontend_tlb_pmp_res_hi_47 = frontend_tlb_pmp__GEN_6 ; 
    wire frontend_tlb_pmp_res_cur_7_cfg_r = frontend_tlb_pmp_io_pmp_0_cfg_r | frontend_tlb_pmp_res_ignore_7 ; 
    wire frontend_tlb_pmp_res_cur_7_cfg_w = frontend_tlb_pmp_io_pmp_0_cfg_w | frontend_tlb_pmp_res_ignore_7 ; 
    wire frontend_tlb_pmp_res_cur_7_cfg_x = frontend_tlb_pmp_io_pmp_0_cfg_x | frontend_tlb_pmp_res_ignore_7 ; 
    wire frontend_tlb_pmp_res_cfg_l = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_l : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_l : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_l : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_l : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_l : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_l : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_l : frontend_tlb_pmp_res_hit & frontend_tlb_pmp_res_cur_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cfg_a = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_a : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_a : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_a : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_a : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_a : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_a : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_a : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_a :2'h0; 
    wire frontend_tlb_pmp_res_cfg_x = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_x : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_x : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_x : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_x : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_x : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_x : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_x : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_x : frontend_tlb_pmp_pmp0_cfg_x ; 
    wire frontend_tlb_pmp_res_cfg_w = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_w : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_w : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_w : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_w : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_w : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_w : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_w : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_w : frontend_tlb_pmp_pmp0_cfg_w ; 
    wire frontend_tlb_pmp_res_cfg_r = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_r : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_r : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_r : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_r : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_r : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_r : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_r : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_r : frontend_tlb_pmp_pmp0_cfg_r ; 
    wire[29:0] frontend_tlb_pmp_res_addr = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_addr : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_addr : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_addr : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_addr : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_addr : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_addr : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_addr : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_addr :30'h0; 
    wire[31:0] frontend_tlb_pmp_res_mask = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_mask : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_mask : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_mask : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_mask : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_mask : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_mask : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_mask : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_mask :32'h0; 
  assign  frontend_tlb_pmp_io_r = frontend_tlb_pmp_res_cfg_r ; 
  assign  frontend_tlb_pmp_io_w = frontend_tlb_pmp_res_cfg_w ; 
  assign  frontend_tlb_pmp_io_x = frontend_tlb_pmp_res_cfg_x ;
    assign frontend_tlb_pmp_io_prv = frontend_tlb_mpu_priv[1:0];
    assign frontend_tlb_pmp_io_pmp_0_cfg_l = frontend_tlb_io_ptw_pmp_0_cfg_l;
    assign frontend_tlb_pmp_io_pmp_0_cfg_a = frontend_tlb_io_ptw_pmp_0_cfg_a;
    assign frontend_tlb_pmp_io_pmp_0_cfg_x = frontend_tlb_io_ptw_pmp_0_cfg_x;
    assign frontend_tlb_pmp_io_pmp_0_cfg_w = frontend_tlb_io_ptw_pmp_0_cfg_w;
    assign frontend_tlb_pmp_io_pmp_0_cfg_r = frontend_tlb_io_ptw_pmp_0_cfg_r;
    assign frontend_tlb_pmp_io_pmp_0_addr = frontend_tlb_io_ptw_pmp_0_addr;
    assign frontend_tlb_pmp_io_pmp_0_mask = frontend_tlb_io_ptw_pmp_0_mask;
    assign frontend_tlb_pmp_io_pmp_1_cfg_l = frontend_tlb_io_ptw_pmp_1_cfg_l;
    assign frontend_tlb_pmp_io_pmp_1_cfg_a = frontend_tlb_io_ptw_pmp_1_cfg_a;
    assign frontend_tlb_pmp_io_pmp_1_cfg_x = frontend_tlb_io_ptw_pmp_1_cfg_x;
    assign frontend_tlb_pmp_io_pmp_1_cfg_w = frontend_tlb_io_ptw_pmp_1_cfg_w;
    assign frontend_tlb_pmp_io_pmp_1_cfg_r = frontend_tlb_io_ptw_pmp_1_cfg_r;
    assign frontend_tlb_pmp_io_pmp_1_addr = frontend_tlb_io_ptw_pmp_1_addr;
    assign frontend_tlb_pmp_io_pmp_1_mask = frontend_tlb_io_ptw_pmp_1_mask;
    assign frontend_tlb_pmp_io_pmp_2_cfg_l = frontend_tlb_io_ptw_pmp_2_cfg_l;
    assign frontend_tlb_pmp_io_pmp_2_cfg_a = frontend_tlb_io_ptw_pmp_2_cfg_a;
    assign frontend_tlb_pmp_io_pmp_2_cfg_x = frontend_tlb_io_ptw_pmp_2_cfg_x;
    assign frontend_tlb_pmp_io_pmp_2_cfg_w = frontend_tlb_io_ptw_pmp_2_cfg_w;
    assign frontend_tlb_pmp_io_pmp_2_cfg_r = frontend_tlb_io_ptw_pmp_2_cfg_r;
    assign frontend_tlb_pmp_io_pmp_2_addr = frontend_tlb_io_ptw_pmp_2_addr;
    assign frontend_tlb_pmp_io_pmp_2_mask = frontend_tlb_io_ptw_pmp_2_mask;
    assign frontend_tlb_pmp_io_pmp_3_cfg_l = frontend_tlb_io_ptw_pmp_3_cfg_l;
    assign frontend_tlb_pmp_io_pmp_3_cfg_a = frontend_tlb_io_ptw_pmp_3_cfg_a;
    assign frontend_tlb_pmp_io_pmp_3_cfg_x = frontend_tlb_io_ptw_pmp_3_cfg_x;
    assign frontend_tlb_pmp_io_pmp_3_cfg_w = frontend_tlb_io_ptw_pmp_3_cfg_w;
    assign frontend_tlb_pmp_io_pmp_3_cfg_r = frontend_tlb_io_ptw_pmp_3_cfg_r;
    assign frontend_tlb_pmp_io_pmp_3_addr = frontend_tlb_io_ptw_pmp_3_addr;
    assign frontend_tlb_pmp_io_pmp_3_mask = frontend_tlb_io_ptw_pmp_3_mask;
    assign frontend_tlb_pmp_io_pmp_4_cfg_l = frontend_tlb_io_ptw_pmp_4_cfg_l;
    assign frontend_tlb_pmp_io_pmp_4_cfg_a = frontend_tlb_io_ptw_pmp_4_cfg_a;
    assign frontend_tlb_pmp_io_pmp_4_cfg_x = frontend_tlb_io_ptw_pmp_4_cfg_x;
    assign frontend_tlb_pmp_io_pmp_4_cfg_w = frontend_tlb_io_ptw_pmp_4_cfg_w;
    assign frontend_tlb_pmp_io_pmp_4_cfg_r = frontend_tlb_io_ptw_pmp_4_cfg_r;
    assign frontend_tlb_pmp_io_pmp_4_addr = frontend_tlb_io_ptw_pmp_4_addr;
    assign frontend_tlb_pmp_io_pmp_4_mask = frontend_tlb_io_ptw_pmp_4_mask;
    assign frontend_tlb_pmp_io_pmp_5_cfg_l = frontend_tlb_io_ptw_pmp_5_cfg_l;
    assign frontend_tlb_pmp_io_pmp_5_cfg_a = frontend_tlb_io_ptw_pmp_5_cfg_a;
    assign frontend_tlb_pmp_io_pmp_5_cfg_x = frontend_tlb_io_ptw_pmp_5_cfg_x;
    assign frontend_tlb_pmp_io_pmp_5_cfg_w = frontend_tlb_io_ptw_pmp_5_cfg_w;
    assign frontend_tlb_pmp_io_pmp_5_cfg_r = frontend_tlb_io_ptw_pmp_5_cfg_r;
    assign frontend_tlb_pmp_io_pmp_5_addr = frontend_tlb_io_ptw_pmp_5_addr;
    assign frontend_tlb_pmp_io_pmp_5_mask = frontend_tlb_io_ptw_pmp_5_mask;
    assign frontend_tlb_pmp_io_pmp_6_cfg_l = frontend_tlb_io_ptw_pmp_6_cfg_l;
    assign frontend_tlb_pmp_io_pmp_6_cfg_a = frontend_tlb_io_ptw_pmp_6_cfg_a;
    assign frontend_tlb_pmp_io_pmp_6_cfg_x = frontend_tlb_io_ptw_pmp_6_cfg_x;
    assign frontend_tlb_pmp_io_pmp_6_cfg_w = frontend_tlb_io_ptw_pmp_6_cfg_w;
    assign frontend_tlb_pmp_io_pmp_6_cfg_r = frontend_tlb_io_ptw_pmp_6_cfg_r;
    assign frontend_tlb_pmp_io_pmp_6_addr = frontend_tlb_io_ptw_pmp_6_addr;
    assign frontend_tlb_pmp_io_pmp_6_mask = frontend_tlb_io_ptw_pmp_6_mask;
    assign frontend_tlb_pmp_io_pmp_7_cfg_l = frontend_tlb_io_ptw_pmp_7_cfg_l;
    assign frontend_tlb_pmp_io_pmp_7_cfg_a = frontend_tlb_io_ptw_pmp_7_cfg_a;
    assign frontend_tlb_pmp_io_pmp_7_cfg_x = frontend_tlb_io_ptw_pmp_7_cfg_x;
    assign frontend_tlb_pmp_io_pmp_7_cfg_w = frontend_tlb_io_ptw_pmp_7_cfg_w;
    assign frontend_tlb_pmp_io_pmp_7_cfg_r = frontend_tlb_io_ptw_pmp_7_cfg_r;
    assign frontend_tlb_pmp_io_pmp_7_addr = frontend_tlb_io_ptw_pmp_7_addr;
    assign frontend_tlb_pmp_io_pmp_7_mask = frontend_tlb_io_ptw_pmp_7_mask;
    assign frontend_tlb_pmp_io_addr = frontend_tlb_mpu_physaddr;
    assign frontend_tlb__pmp_io_r = frontend_tlb_pmp_io_r;
    assign frontend_tlb__pmp_io_w = frontend_tlb_pmp_io_w;
    assign frontend_tlb__pmp_io_x = frontend_tlb_pmp_io_x;
      
    wire frontend_tlb_entries_barrier_io_x_u;
    wire frontend_tlb_entries_barrier_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_io_x_ae_final;
    wire frontend_tlb_entries_barrier_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_io_x_pf;
    wire frontend_tlb_entries_barrier_io_x_gf;
    wire frontend_tlb_entries_barrier_io_x_sw;
    wire frontend_tlb_entries_barrier_io_x_sx;
    wire frontend_tlb_entries_barrier_io_x_sr;
    wire frontend_tlb_entries_barrier_io_x_hw;
    wire frontend_tlb_entries_barrier_io_x_hx;
    wire frontend_tlb_entries_barrier_io_x_hr;
    wire frontend_tlb_entries_barrier_io_x_pw;
    wire frontend_tlb_entries_barrier_io_x_px;
    wire frontend_tlb_entries_barrier_io_x_pr;
    wire frontend_tlb_entries_barrier_io_x_ppp;
    wire frontend_tlb_entries_barrier_io_x_pal;
    wire frontend_tlb_entries_barrier_io_x_paa;
    wire frontend_tlb_entries_barrier_io_x_eff;
    wire frontend_tlb_entries_barrier_io_x_c;
    wire frontend_tlb_entries_barrier_io_y_u;
    wire frontend_tlb_entries_barrier_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_io_y_ae_final;
    wire frontend_tlb_entries_barrier_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_io_y_pf;
    wire frontend_tlb_entries_barrier_io_y_gf;
    wire frontend_tlb_entries_barrier_io_y_sw;
    wire frontend_tlb_entries_barrier_io_y_sx;
    wire frontend_tlb_entries_barrier_io_y_sr;
    wire frontend_tlb_entries_barrier_io_y_hw;
    wire frontend_tlb_entries_barrier_io_y_hx;
    wire frontend_tlb_entries_barrier_io_y_hr;
    wire frontend_tlb_entries_barrier_io_y_pw;
    wire frontend_tlb_entries_barrier_io_y_px;
    wire frontend_tlb_entries_barrier_io_y_pr;
    wire frontend_tlb_entries_barrier_io_y_ppp;
    wire frontend_tlb_entries_barrier_io_y_pal;
    wire frontend_tlb_entries_barrier_io_y_paa;
    wire frontend_tlb_entries_barrier_io_y_eff;
    wire frontend_tlb_entries_barrier_io_y_c;
    wire frontend_tlb_entries_barrier_1_io_x_u;
    wire frontend_tlb_entries_barrier_1_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_1_io_x_ae_final;
    wire frontend_tlb_entries_barrier_1_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_1_io_x_pf;
    wire frontend_tlb_entries_barrier_1_io_x_gf;
    wire frontend_tlb_entries_barrier_1_io_x_sw;
    wire frontend_tlb_entries_barrier_1_io_x_sx;
    wire frontend_tlb_entries_barrier_1_io_x_sr;
    wire frontend_tlb_entries_barrier_1_io_x_hw;
    wire frontend_tlb_entries_barrier_1_io_x_hx;
    wire frontend_tlb_entries_barrier_1_io_x_hr;
    wire frontend_tlb_entries_barrier_1_io_x_pw;
    wire frontend_tlb_entries_barrier_1_io_x_px;
    wire frontend_tlb_entries_barrier_1_io_x_pr;
    wire frontend_tlb_entries_barrier_1_io_x_ppp;
    wire frontend_tlb_entries_barrier_1_io_x_pal;
    wire frontend_tlb_entries_barrier_1_io_x_paa;
    wire frontend_tlb_entries_barrier_1_io_x_eff;
    wire frontend_tlb_entries_barrier_1_io_x_c;
    wire frontend_tlb_entries_barrier_1_io_y_u;
    wire frontend_tlb_entries_barrier_1_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_1_io_y_ae_final;
    wire frontend_tlb_entries_barrier_1_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_1_io_y_pf;
    wire frontend_tlb_entries_barrier_1_io_y_gf;
    wire frontend_tlb_entries_barrier_1_io_y_sw;
    wire frontend_tlb_entries_barrier_1_io_y_sx;
    wire frontend_tlb_entries_barrier_1_io_y_sr;
    wire frontend_tlb_entries_barrier_1_io_y_hw;
    wire frontend_tlb_entries_barrier_1_io_y_hx;
    wire frontend_tlb_entries_barrier_1_io_y_hr;
    wire frontend_tlb_entries_barrier_1_io_y_pw;
    wire frontend_tlb_entries_barrier_1_io_y_px;
    wire frontend_tlb_entries_barrier_1_io_y_pr;
    wire frontend_tlb_entries_barrier_1_io_y_ppp;
    wire frontend_tlb_entries_barrier_1_io_y_pal;
    wire frontend_tlb_entries_barrier_1_io_y_paa;
    wire frontend_tlb_entries_barrier_1_io_y_eff;
    wire frontend_tlb_entries_barrier_1_io_y_c;
    wire frontend_tlb_entries_barrier_2_io_x_u;
    wire frontend_tlb_entries_barrier_2_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_2_io_x_ae_final;
    wire frontend_tlb_entries_barrier_2_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_2_io_x_pf;
    wire frontend_tlb_entries_barrier_2_io_x_gf;
    wire frontend_tlb_entries_barrier_2_io_x_sw;
    wire frontend_tlb_entries_barrier_2_io_x_sx;
    wire frontend_tlb_entries_barrier_2_io_x_sr;
    wire frontend_tlb_entries_barrier_2_io_x_hw;
    wire frontend_tlb_entries_barrier_2_io_x_hx;
    wire frontend_tlb_entries_barrier_2_io_x_hr;
    wire frontend_tlb_entries_barrier_2_io_x_pw;
    wire frontend_tlb_entries_barrier_2_io_x_px;
    wire frontend_tlb_entries_barrier_2_io_x_pr;
    wire frontend_tlb_entries_barrier_2_io_x_ppp;
    wire frontend_tlb_entries_barrier_2_io_x_pal;
    wire frontend_tlb_entries_barrier_2_io_x_paa;
    wire frontend_tlb_entries_barrier_2_io_x_eff;
    wire frontend_tlb_entries_barrier_2_io_x_c;
    wire frontend_tlb_entries_barrier_2_io_y_u;
    wire frontend_tlb_entries_barrier_2_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_2_io_y_ae_final;
    wire frontend_tlb_entries_barrier_2_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_2_io_y_pf;
    wire frontend_tlb_entries_barrier_2_io_y_gf;
    wire frontend_tlb_entries_barrier_2_io_y_sw;
    wire frontend_tlb_entries_barrier_2_io_y_sx;
    wire frontend_tlb_entries_barrier_2_io_y_sr;
    wire frontend_tlb_entries_barrier_2_io_y_hw;
    wire frontend_tlb_entries_barrier_2_io_y_hx;
    wire frontend_tlb_entries_barrier_2_io_y_hr;
    wire frontend_tlb_entries_barrier_2_io_y_pw;
    wire frontend_tlb_entries_barrier_2_io_y_px;
    wire frontend_tlb_entries_barrier_2_io_y_pr;
    wire frontend_tlb_entries_barrier_2_io_y_ppp;
    wire frontend_tlb_entries_barrier_2_io_y_pal;
    wire frontend_tlb_entries_barrier_2_io_y_paa;
    wire frontend_tlb_entries_barrier_2_io_y_eff;
    wire frontend_tlb_entries_barrier_2_io_y_c;
    wire frontend_tlb_entries_barrier_3_io_x_u;
    wire frontend_tlb_entries_barrier_3_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_3_io_x_ae_final;
    wire frontend_tlb_entries_barrier_3_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_3_io_x_pf;
    wire frontend_tlb_entries_barrier_3_io_x_gf;
    wire frontend_tlb_entries_barrier_3_io_x_sw;
    wire frontend_tlb_entries_barrier_3_io_x_sx;
    wire frontend_tlb_entries_barrier_3_io_x_sr;
    wire frontend_tlb_entries_barrier_3_io_x_hw;
    wire frontend_tlb_entries_barrier_3_io_x_hx;
    wire frontend_tlb_entries_barrier_3_io_x_hr;
    wire frontend_tlb_entries_barrier_3_io_x_pw;
    wire frontend_tlb_entries_barrier_3_io_x_px;
    wire frontend_tlb_entries_barrier_3_io_x_pr;
    wire frontend_tlb_entries_barrier_3_io_x_ppp;
    wire frontend_tlb_entries_barrier_3_io_x_pal;
    wire frontend_tlb_entries_barrier_3_io_x_paa;
    wire frontend_tlb_entries_barrier_3_io_x_eff;
    wire frontend_tlb_entries_barrier_3_io_x_c;
    wire frontend_tlb_entries_barrier_3_io_y_u;
    wire frontend_tlb_entries_barrier_3_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_3_io_y_ae_final;
    wire frontend_tlb_entries_barrier_3_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_3_io_y_pf;
    wire frontend_tlb_entries_barrier_3_io_y_gf;
    wire frontend_tlb_entries_barrier_3_io_y_sw;
    wire frontend_tlb_entries_barrier_3_io_y_sx;
    wire frontend_tlb_entries_barrier_3_io_y_sr;
    wire frontend_tlb_entries_barrier_3_io_y_hw;
    wire frontend_tlb_entries_barrier_3_io_y_hx;
    wire frontend_tlb_entries_barrier_3_io_y_hr;
    wire frontend_tlb_entries_barrier_3_io_y_pw;
    wire frontend_tlb_entries_barrier_3_io_y_px;
    wire frontend_tlb_entries_barrier_3_io_y_pr;
    wire frontend_tlb_entries_barrier_3_io_y_ppp;
    wire frontend_tlb_entries_barrier_3_io_y_pal;
    wire frontend_tlb_entries_barrier_3_io_y_paa;
    wire frontend_tlb_entries_barrier_3_io_y_eff;
    wire frontend_tlb_entries_barrier_3_io_y_c;
    wire frontend_tlb_entries_barrier_4_io_x_u;
    wire frontend_tlb_entries_barrier_4_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_4_io_x_ae_final;
    wire frontend_tlb_entries_barrier_4_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_4_io_x_pf;
    wire frontend_tlb_entries_barrier_4_io_x_gf;
    wire frontend_tlb_entries_barrier_4_io_x_sw;
    wire frontend_tlb_entries_barrier_4_io_x_sx;
    wire frontend_tlb_entries_barrier_4_io_x_sr;
    wire frontend_tlb_entries_barrier_4_io_x_hw;
    wire frontend_tlb_entries_barrier_4_io_x_hx;
    wire frontend_tlb_entries_barrier_4_io_x_hr;
    wire frontend_tlb_entries_barrier_4_io_x_pw;
    wire frontend_tlb_entries_barrier_4_io_x_px;
    wire frontend_tlb_entries_barrier_4_io_x_pr;
    wire frontend_tlb_entries_barrier_4_io_x_ppp;
    wire frontend_tlb_entries_barrier_4_io_x_pal;
    wire frontend_tlb_entries_barrier_4_io_x_paa;
    wire frontend_tlb_entries_barrier_4_io_x_eff;
    wire frontend_tlb_entries_barrier_4_io_x_c;
    wire frontend_tlb_entries_barrier_4_io_y_u;
    wire frontend_tlb_entries_barrier_4_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_4_io_y_ae_final;
    wire frontend_tlb_entries_barrier_4_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_4_io_y_pf;
    wire frontend_tlb_entries_barrier_4_io_y_gf;
    wire frontend_tlb_entries_barrier_4_io_y_sw;
    wire frontend_tlb_entries_barrier_4_io_y_sx;
    wire frontend_tlb_entries_barrier_4_io_y_sr;
    wire frontend_tlb_entries_barrier_4_io_y_hw;
    wire frontend_tlb_entries_barrier_4_io_y_hx;
    wire frontend_tlb_entries_barrier_4_io_y_hr;
    wire frontend_tlb_entries_barrier_4_io_y_pw;
    wire frontend_tlb_entries_barrier_4_io_y_px;
    wire frontend_tlb_entries_barrier_4_io_y_pr;
    wire frontend_tlb_entries_barrier_4_io_y_ppp;
    wire frontend_tlb_entries_barrier_4_io_y_pal;
    wire frontend_tlb_entries_barrier_4_io_y_paa;
    wire frontend_tlb_entries_barrier_4_io_y_eff;
    wire frontend_tlb_entries_barrier_4_io_y_c;
    wire frontend_tlb_entries_barrier_5_io_x_u;
    wire frontend_tlb_entries_barrier_5_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_5_io_x_ae_final;
    wire frontend_tlb_entries_barrier_5_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_5_io_x_pf;
    wire frontend_tlb_entries_barrier_5_io_x_gf;
    wire frontend_tlb_entries_barrier_5_io_x_sw;
    wire frontend_tlb_entries_barrier_5_io_x_sx;
    wire frontend_tlb_entries_barrier_5_io_x_sr;
    wire frontend_tlb_entries_barrier_5_io_x_hw;
    wire frontend_tlb_entries_barrier_5_io_x_hx;
    wire frontend_tlb_entries_barrier_5_io_x_hr;
    wire frontend_tlb_entries_barrier_5_io_x_pw;
    wire frontend_tlb_entries_barrier_5_io_x_px;
    wire frontend_tlb_entries_barrier_5_io_x_pr;
    wire frontend_tlb_entries_barrier_5_io_x_ppp;
    wire frontend_tlb_entries_barrier_5_io_x_pal;
    wire frontend_tlb_entries_barrier_5_io_x_paa;
    wire frontend_tlb_entries_barrier_5_io_x_eff;
    wire frontend_tlb_entries_barrier_5_io_x_c;
    wire frontend_tlb_entries_barrier_5_io_y_u;
    wire frontend_tlb_entries_barrier_5_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_5_io_y_ae_final;
    wire frontend_tlb_entries_barrier_5_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_5_io_y_pf;
    wire frontend_tlb_entries_barrier_5_io_y_gf;
    wire frontend_tlb_entries_barrier_5_io_y_sw;
    wire frontend_tlb_entries_barrier_5_io_y_sx;
    wire frontend_tlb_entries_barrier_5_io_y_sr;
    wire frontend_tlb_entries_barrier_5_io_y_hw;
    wire frontend_tlb_entries_barrier_5_io_y_hx;
    wire frontend_tlb_entries_barrier_5_io_y_hr;
    wire frontend_tlb_entries_barrier_5_io_y_pw;
    wire frontend_tlb_entries_barrier_5_io_y_px;
    wire frontend_tlb_entries_barrier_5_io_y_pr;
    wire frontend_tlb_entries_barrier_5_io_y_ppp;
    wire frontend_tlb_entries_barrier_5_io_y_pal;
    wire frontend_tlb_entries_barrier_5_io_y_paa;
    wire frontend_tlb_entries_barrier_5_io_y_eff;
    wire frontend_tlb_entries_barrier_5_io_y_c;

    assign  frontend_tlb_entries_barrier_io_y_u = frontend_tlb_entries_barrier_io_x_u ; 
  assign  frontend_tlb_entries_barrier_io_y_ae_ptw = frontend_tlb_entries_barrier_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_io_y_ae_final = frontend_tlb_entries_barrier_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_io_y_ae_stage2 = frontend_tlb_entries_barrier_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_io_y_pf = frontend_tlb_entries_barrier_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_io_y_gf = frontend_tlb_entries_barrier_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_io_y_sw = frontend_tlb_entries_barrier_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_io_y_sx = frontend_tlb_entries_barrier_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_io_y_sr = frontend_tlb_entries_barrier_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_io_y_hw = frontend_tlb_entries_barrier_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_io_y_hx = frontend_tlb_entries_barrier_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_io_y_hr = frontend_tlb_entries_barrier_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_io_y_pw = frontend_tlb_entries_barrier_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_io_y_px = frontend_tlb_entries_barrier_io_x_px ; 
  assign  frontend_tlb_entries_barrier_io_y_pr = frontend_tlb_entries_barrier_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_io_y_ppp = frontend_tlb_entries_barrier_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_io_y_pal = frontend_tlb_entries_barrier_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_io_y_paa = frontend_tlb_entries_barrier_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_io_y_eff = frontend_tlb_entries_barrier_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_io_y_c = frontend_tlb_entries_barrier_io_x_c ;
    assign  frontend_tlb_entries_barrier_1_io_y_u = frontend_tlb_entries_barrier_1_io_x_u ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ae_ptw = frontend_tlb_entries_barrier_1_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ae_final = frontend_tlb_entries_barrier_1_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ae_stage2 = frontend_tlb_entries_barrier_1_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pf = frontend_tlb_entries_barrier_1_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_1_io_y_gf = frontend_tlb_entries_barrier_1_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_1_io_y_sw = frontend_tlb_entries_barrier_1_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_sx = frontend_tlb_entries_barrier_1_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_1_io_y_sr = frontend_tlb_entries_barrier_1_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_1_io_y_hw = frontend_tlb_entries_barrier_1_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_hx = frontend_tlb_entries_barrier_1_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_1_io_y_hr = frontend_tlb_entries_barrier_1_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pw = frontend_tlb_entries_barrier_1_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_px = frontend_tlb_entries_barrier_1_io_x_px ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pr = frontend_tlb_entries_barrier_1_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ppp = frontend_tlb_entries_barrier_1_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pal = frontend_tlb_entries_barrier_1_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_1_io_y_paa = frontend_tlb_entries_barrier_1_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_1_io_y_eff = frontend_tlb_entries_barrier_1_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_1_io_y_c = frontend_tlb_entries_barrier_1_io_x_c ;
    assign  frontend_tlb_entries_barrier_2_io_y_u = frontend_tlb_entries_barrier_2_io_x_u ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ae_ptw = frontend_tlb_entries_barrier_2_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ae_final = frontend_tlb_entries_barrier_2_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ae_stage2 = frontend_tlb_entries_barrier_2_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pf = frontend_tlb_entries_barrier_2_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_2_io_y_gf = frontend_tlb_entries_barrier_2_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_2_io_y_sw = frontend_tlb_entries_barrier_2_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_sx = frontend_tlb_entries_barrier_2_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_2_io_y_sr = frontend_tlb_entries_barrier_2_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_2_io_y_hw = frontend_tlb_entries_barrier_2_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_hx = frontend_tlb_entries_barrier_2_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_2_io_y_hr = frontend_tlb_entries_barrier_2_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pw = frontend_tlb_entries_barrier_2_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_px = frontend_tlb_entries_barrier_2_io_x_px ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pr = frontend_tlb_entries_barrier_2_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ppp = frontend_tlb_entries_barrier_2_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pal = frontend_tlb_entries_barrier_2_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_2_io_y_paa = frontend_tlb_entries_barrier_2_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_2_io_y_eff = frontend_tlb_entries_barrier_2_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_2_io_y_c = frontend_tlb_entries_barrier_2_io_x_c ;
    assign  frontend_tlb_entries_barrier_3_io_y_u = frontend_tlb_entries_barrier_3_io_x_u ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ae_ptw = frontend_tlb_entries_barrier_3_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ae_final = frontend_tlb_entries_barrier_3_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ae_stage2 = frontend_tlb_entries_barrier_3_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pf = frontend_tlb_entries_barrier_3_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_3_io_y_gf = frontend_tlb_entries_barrier_3_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_3_io_y_sw = frontend_tlb_entries_barrier_3_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_sx = frontend_tlb_entries_barrier_3_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_3_io_y_sr = frontend_tlb_entries_barrier_3_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_3_io_y_hw = frontend_tlb_entries_barrier_3_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_hx = frontend_tlb_entries_barrier_3_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_3_io_y_hr = frontend_tlb_entries_barrier_3_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pw = frontend_tlb_entries_barrier_3_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_px = frontend_tlb_entries_barrier_3_io_x_px ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pr = frontend_tlb_entries_barrier_3_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ppp = frontend_tlb_entries_barrier_3_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pal = frontend_tlb_entries_barrier_3_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_3_io_y_paa = frontend_tlb_entries_barrier_3_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_3_io_y_eff = frontend_tlb_entries_barrier_3_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_3_io_y_c = frontend_tlb_entries_barrier_3_io_x_c ;
    assign  frontend_tlb_entries_barrier_4_io_y_u = frontend_tlb_entries_barrier_4_io_x_u ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ae_ptw = frontend_tlb_entries_barrier_4_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ae_final = frontend_tlb_entries_barrier_4_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ae_stage2 = frontend_tlb_entries_barrier_4_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pf = frontend_tlb_entries_barrier_4_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_4_io_y_gf = frontend_tlb_entries_barrier_4_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_4_io_y_sw = frontend_tlb_entries_barrier_4_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_sx = frontend_tlb_entries_barrier_4_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_4_io_y_sr = frontend_tlb_entries_barrier_4_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_4_io_y_hw = frontend_tlb_entries_barrier_4_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_hx = frontend_tlb_entries_barrier_4_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_4_io_y_hr = frontend_tlb_entries_barrier_4_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pw = frontend_tlb_entries_barrier_4_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_px = frontend_tlb_entries_barrier_4_io_x_px ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pr = frontend_tlb_entries_barrier_4_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ppp = frontend_tlb_entries_barrier_4_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pal = frontend_tlb_entries_barrier_4_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_4_io_y_paa = frontend_tlb_entries_barrier_4_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_4_io_y_eff = frontend_tlb_entries_barrier_4_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_4_io_y_c = frontend_tlb_entries_barrier_4_io_x_c ;
    assign  frontend_tlb_entries_barrier_5_io_y_u = frontend_tlb_entries_barrier_5_io_x_u ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ae_ptw = frontend_tlb_entries_barrier_5_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ae_final = frontend_tlb_entries_barrier_5_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ae_stage2 = frontend_tlb_entries_barrier_5_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pf = frontend_tlb_entries_barrier_5_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_5_io_y_gf = frontend_tlb_entries_barrier_5_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_5_io_y_sw = frontend_tlb_entries_barrier_5_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_sx = frontend_tlb_entries_barrier_5_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_5_io_y_sr = frontend_tlb_entries_barrier_5_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_5_io_y_hw = frontend_tlb_entries_barrier_5_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_hx = frontend_tlb_entries_barrier_5_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_5_io_y_hr = frontend_tlb_entries_barrier_5_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pw = frontend_tlb_entries_barrier_5_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_px = frontend_tlb_entries_barrier_5_io_x_px ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pr = frontend_tlb_entries_barrier_5_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ppp = frontend_tlb_entries_barrier_5_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pal = frontend_tlb_entries_barrier_5_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_5_io_y_paa = frontend_tlb_entries_barrier_5_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_5_io_y_eff = frontend_tlb_entries_barrier_5_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_5_io_y_c = frontend_tlb_entries_barrier_5_io_x_c ;
    assign frontend_tlb_entries_barrier_io_x_u = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_ae_ptw = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_ae_final = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_ae_stage2 = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_pf = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_gf = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_sw = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_sx = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_sr = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_hw = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_hx = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_hr = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_pw = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_px = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_pr = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_ppp = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_pal = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_paa = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_eff = 1'h0;
    assign frontend_tlb_entries_barrier_io_x_c = 1'h0;
    assign frontend_tlb__entries_barrier_io_y_u = frontend_tlb_entries_barrier_io_y_u;
    assign frontend_tlb__entries_barrier_io_y_ae_ptw = frontend_tlb_entries_barrier_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_io_y_ae_final = frontend_tlb_entries_barrier_io_y_ae_final;
    assign frontend_tlb__entries_barrier_io_y_ae_stage2 = frontend_tlb_entries_barrier_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_io_y_pf = frontend_tlb_entries_barrier_io_y_pf;
    assign frontend_tlb__entries_barrier_io_y_gf = frontend_tlb_entries_barrier_io_y_gf;
    assign frontend_tlb__entries_barrier_io_y_sw = frontend_tlb_entries_barrier_io_y_sw;
    assign frontend_tlb__entries_barrier_io_y_sx = frontend_tlb_entries_barrier_io_y_sx;
    assign frontend_tlb__entries_barrier_io_y_sr = frontend_tlb_entries_barrier_io_y_sr;
    assign frontend_tlb__entries_barrier_io_y_hw = frontend_tlb_entries_barrier_io_y_hw;
    assign frontend_tlb__entries_barrier_io_y_hx = frontend_tlb_entries_barrier_io_y_hx;
    assign frontend_tlb__entries_barrier_io_y_hr = frontend_tlb_entries_barrier_io_y_hr;
    assign frontend_tlb__entries_barrier_io_y_pw = frontend_tlb_entries_barrier_io_y_pw;
    assign frontend_tlb__entries_barrier_io_y_px = frontend_tlb_entries_barrier_io_y_px;
    assign frontend_tlb__entries_barrier_io_y_pr = frontend_tlb_entries_barrier_io_y_pr;
    assign frontend_tlb__entries_barrier_io_y_ppp = frontend_tlb_entries_barrier_io_y_ppp;
    assign frontend_tlb__entries_barrier_io_y_pal = frontend_tlb_entries_barrier_io_y_pal;
    assign frontend_tlb__entries_barrier_io_y_paa = frontend_tlb_entries_barrier_io_y_paa;
    assign frontend_tlb__entries_barrier_io_y_eff = frontend_tlb_entries_barrier_io_y_eff;
    assign frontend_tlb__entries_barrier_io_y_c = frontend_tlb_entries_barrier_io_y_c;
    assign frontend_tlb_entries_barrier_1_io_x_u = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_ae_ptw = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_ae_final = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_ae_stage2 = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_pf = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_gf = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_sw = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_sx = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_sr = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_hw = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_hx = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_hr = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_pw = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_px = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_pr = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_ppp = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_pal = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_paa = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_eff = 1'h0;
    assign frontend_tlb_entries_barrier_1_io_x_c = 1'h0;
    assign frontend_tlb__entries_barrier_1_io_y_u = frontend_tlb_entries_barrier_1_io_y_u;
    assign frontend_tlb__entries_barrier_1_io_y_ae_ptw = frontend_tlb_entries_barrier_1_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_1_io_y_ae_final = frontend_tlb_entries_barrier_1_io_y_ae_final;
    assign frontend_tlb__entries_barrier_1_io_y_ae_stage2 = frontend_tlb_entries_barrier_1_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_1_io_y_pf = frontend_tlb_entries_barrier_1_io_y_pf;
    assign frontend_tlb__entries_barrier_1_io_y_gf = frontend_tlb_entries_barrier_1_io_y_gf;
    assign frontend_tlb__entries_barrier_1_io_y_sw = frontend_tlb_entries_barrier_1_io_y_sw;
    assign frontend_tlb__entries_barrier_1_io_y_sx = frontend_tlb_entries_barrier_1_io_y_sx;
    assign frontend_tlb__entries_barrier_1_io_y_sr = frontend_tlb_entries_barrier_1_io_y_sr;
    assign frontend_tlb__entries_barrier_1_io_y_hw = frontend_tlb_entries_barrier_1_io_y_hw;
    assign frontend_tlb__entries_barrier_1_io_y_hx = frontend_tlb_entries_barrier_1_io_y_hx;
    assign frontend_tlb__entries_barrier_1_io_y_hr = frontend_tlb_entries_barrier_1_io_y_hr;
    assign frontend_tlb__entries_barrier_1_io_y_pw = frontend_tlb_entries_barrier_1_io_y_pw;
    assign frontend_tlb__entries_barrier_1_io_y_px = frontend_tlb_entries_barrier_1_io_y_px;
    assign frontend_tlb__entries_barrier_1_io_y_pr = frontend_tlb_entries_barrier_1_io_y_pr;
    assign frontend_tlb__entries_barrier_1_io_y_ppp = frontend_tlb_entries_barrier_1_io_y_ppp;
    assign frontend_tlb__entries_barrier_1_io_y_pal = frontend_tlb_entries_barrier_1_io_y_pal;
    assign frontend_tlb__entries_barrier_1_io_y_paa = frontend_tlb_entries_barrier_1_io_y_paa;
    assign frontend_tlb__entries_barrier_1_io_y_eff = frontend_tlb_entries_barrier_1_io_y_eff;
    assign frontend_tlb__entries_barrier_1_io_y_c = frontend_tlb_entries_barrier_1_io_y_c;
    assign frontend_tlb_entries_barrier_2_io_x_u = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_ae_ptw = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_ae_final = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_ae_stage2 = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_pf = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_gf = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_sw = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_sx = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_sr = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_hw = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_hx = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_hr = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_pw = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_px = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_pr = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_ppp = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_pal = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_paa = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_eff = 1'h0;
    assign frontend_tlb_entries_barrier_2_io_x_c = 1'h0;
    assign frontend_tlb__entries_barrier_2_io_y_u = frontend_tlb_entries_barrier_2_io_y_u;
    assign frontend_tlb__entries_barrier_2_io_y_ae_ptw = frontend_tlb_entries_barrier_2_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_2_io_y_ae_final = frontend_tlb_entries_barrier_2_io_y_ae_final;
    assign frontend_tlb__entries_barrier_2_io_y_ae_stage2 = frontend_tlb_entries_barrier_2_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_2_io_y_pf = frontend_tlb_entries_barrier_2_io_y_pf;
    assign frontend_tlb__entries_barrier_2_io_y_gf = frontend_tlb_entries_barrier_2_io_y_gf;
    assign frontend_tlb__entries_barrier_2_io_y_sw = frontend_tlb_entries_barrier_2_io_y_sw;
    assign frontend_tlb__entries_barrier_2_io_y_sx = frontend_tlb_entries_barrier_2_io_y_sx;
    assign frontend_tlb__entries_barrier_2_io_y_sr = frontend_tlb_entries_barrier_2_io_y_sr;
    assign frontend_tlb__entries_barrier_2_io_y_hw = frontend_tlb_entries_barrier_2_io_y_hw;
    assign frontend_tlb__entries_barrier_2_io_y_hx = frontend_tlb_entries_barrier_2_io_y_hx;
    assign frontend_tlb__entries_barrier_2_io_y_hr = frontend_tlb_entries_barrier_2_io_y_hr;
    assign frontend_tlb__entries_barrier_2_io_y_pw = frontend_tlb_entries_barrier_2_io_y_pw;
    assign frontend_tlb__entries_barrier_2_io_y_px = frontend_tlb_entries_barrier_2_io_y_px;
    assign frontend_tlb__entries_barrier_2_io_y_pr = frontend_tlb_entries_barrier_2_io_y_pr;
    assign frontend_tlb__entries_barrier_2_io_y_ppp = frontend_tlb_entries_barrier_2_io_y_ppp;
    assign frontend_tlb__entries_barrier_2_io_y_pal = frontend_tlb_entries_barrier_2_io_y_pal;
    assign frontend_tlb__entries_barrier_2_io_y_paa = frontend_tlb_entries_barrier_2_io_y_paa;
    assign frontend_tlb__entries_barrier_2_io_y_eff = frontend_tlb_entries_barrier_2_io_y_eff;
    assign frontend_tlb__entries_barrier_2_io_y_c = frontend_tlb_entries_barrier_2_io_y_c;
    assign frontend_tlb_entries_barrier_3_io_x_u = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_ae_ptw = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_ae_final = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_ae_stage2 = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_pf = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_gf = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_sw = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_sx = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_sr = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_hw = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_hx = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_hr = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_pw = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_px = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_pr = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_ppp = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_pal = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_paa = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_eff = 1'h0;
    assign frontend_tlb_entries_barrier_3_io_x_c = 1'h0;
    assign frontend_tlb__entries_barrier_3_io_y_u = frontend_tlb_entries_barrier_3_io_y_u;
    assign frontend_tlb__entries_barrier_3_io_y_ae_ptw = frontend_tlb_entries_barrier_3_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_3_io_y_ae_final = frontend_tlb_entries_barrier_3_io_y_ae_final;
    assign frontend_tlb__entries_barrier_3_io_y_ae_stage2 = frontend_tlb_entries_barrier_3_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_3_io_y_pf = frontend_tlb_entries_barrier_3_io_y_pf;
    assign frontend_tlb__entries_barrier_3_io_y_gf = frontend_tlb_entries_barrier_3_io_y_gf;
    assign frontend_tlb__entries_barrier_3_io_y_sw = frontend_tlb_entries_barrier_3_io_y_sw;
    assign frontend_tlb__entries_barrier_3_io_y_sx = frontend_tlb_entries_barrier_3_io_y_sx;
    assign frontend_tlb__entries_barrier_3_io_y_sr = frontend_tlb_entries_barrier_3_io_y_sr;
    assign frontend_tlb__entries_barrier_3_io_y_hw = frontend_tlb_entries_barrier_3_io_y_hw;
    assign frontend_tlb__entries_barrier_3_io_y_hx = frontend_tlb_entries_barrier_3_io_y_hx;
    assign frontend_tlb__entries_barrier_3_io_y_hr = frontend_tlb_entries_barrier_3_io_y_hr;
    assign frontend_tlb__entries_barrier_3_io_y_pw = frontend_tlb_entries_barrier_3_io_y_pw;
    assign frontend_tlb__entries_barrier_3_io_y_px = frontend_tlb_entries_barrier_3_io_y_px;
    assign frontend_tlb__entries_barrier_3_io_y_pr = frontend_tlb_entries_barrier_3_io_y_pr;
    assign frontend_tlb__entries_barrier_3_io_y_ppp = frontend_tlb_entries_barrier_3_io_y_ppp;
    assign frontend_tlb__entries_barrier_3_io_y_pal = frontend_tlb_entries_barrier_3_io_y_pal;
    assign frontend_tlb__entries_barrier_3_io_y_paa = frontend_tlb_entries_barrier_3_io_y_paa;
    assign frontend_tlb__entries_barrier_3_io_y_eff = frontend_tlb_entries_barrier_3_io_y_eff;
    assign frontend_tlb__entries_barrier_3_io_y_c = frontend_tlb_entries_barrier_3_io_y_c;
    assign frontend_tlb_entries_barrier_4_io_x_u = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_ae_ptw = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_ae_final = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_ae_stage2 = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_pf = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_gf = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_sw = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_sx = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_sr = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_hw = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_hx = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_hr = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_pw = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_px = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_pr = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_ppp = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_pal = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_paa = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_eff = 1'h0;
    assign frontend_tlb_entries_barrier_4_io_x_c = 1'h0;
    assign frontend_tlb__entries_barrier_4_io_y_u = frontend_tlb_entries_barrier_4_io_y_u;
    assign frontend_tlb__entries_barrier_4_io_y_ae_ptw = frontend_tlb_entries_barrier_4_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_4_io_y_ae_final = frontend_tlb_entries_barrier_4_io_y_ae_final;
    assign frontend_tlb__entries_barrier_4_io_y_ae_stage2 = frontend_tlb_entries_barrier_4_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_4_io_y_pf = frontend_tlb_entries_barrier_4_io_y_pf;
    assign frontend_tlb__entries_barrier_4_io_y_gf = frontend_tlb_entries_barrier_4_io_y_gf;
    assign frontend_tlb__entries_barrier_4_io_y_sw = frontend_tlb_entries_barrier_4_io_y_sw;
    assign frontend_tlb__entries_barrier_4_io_y_sx = frontend_tlb_entries_barrier_4_io_y_sx;
    assign frontend_tlb__entries_barrier_4_io_y_sr = frontend_tlb_entries_barrier_4_io_y_sr;
    assign frontend_tlb__entries_barrier_4_io_y_hw = frontend_tlb_entries_barrier_4_io_y_hw;
    assign frontend_tlb__entries_barrier_4_io_y_hx = frontend_tlb_entries_barrier_4_io_y_hx;
    assign frontend_tlb__entries_barrier_4_io_y_hr = frontend_tlb_entries_barrier_4_io_y_hr;
    assign frontend_tlb__entries_barrier_4_io_y_pw = frontend_tlb_entries_barrier_4_io_y_pw;
    assign frontend_tlb__entries_barrier_4_io_y_px = frontend_tlb_entries_barrier_4_io_y_px;
    assign frontend_tlb__entries_barrier_4_io_y_pr = frontend_tlb_entries_barrier_4_io_y_pr;
    assign frontend_tlb__entries_barrier_4_io_y_ppp = frontend_tlb_entries_barrier_4_io_y_ppp;
    assign frontend_tlb__entries_barrier_4_io_y_pal = frontend_tlb_entries_barrier_4_io_y_pal;
    assign frontend_tlb__entries_barrier_4_io_y_paa = frontend_tlb_entries_barrier_4_io_y_paa;
    assign frontend_tlb__entries_barrier_4_io_y_eff = frontend_tlb_entries_barrier_4_io_y_eff;
    assign frontend_tlb__entries_barrier_4_io_y_c = frontend_tlb_entries_barrier_4_io_y_c;
    assign frontend_tlb_entries_barrier_5_io_x_u = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_ae_ptw = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_ae_final = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_ae_stage2 = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_pf = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_gf = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_sw = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_sx = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_sr = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_hw = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_hx = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_hr = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_pw = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_px = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_pr = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_ppp = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_pal = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_paa = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_eff = 1'h0;
    assign frontend_tlb_entries_barrier_5_io_x_c = 1'h0;
    assign frontend_tlb__entries_barrier_5_io_y_u = frontend_tlb_entries_barrier_5_io_y_u;
    assign frontend_tlb__entries_barrier_5_io_y_ae_ptw = frontend_tlb_entries_barrier_5_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_5_io_y_ae_final = frontend_tlb_entries_barrier_5_io_y_ae_final;
    assign frontend_tlb__entries_barrier_5_io_y_ae_stage2 = frontend_tlb_entries_barrier_5_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_5_io_y_pf = frontend_tlb_entries_barrier_5_io_y_pf;
    assign frontend_tlb__entries_barrier_5_io_y_gf = frontend_tlb_entries_barrier_5_io_y_gf;
    assign frontend_tlb__entries_barrier_5_io_y_sw = frontend_tlb_entries_barrier_5_io_y_sw;
    assign frontend_tlb__entries_barrier_5_io_y_sx = frontend_tlb_entries_barrier_5_io_y_sx;
    assign frontend_tlb__entries_barrier_5_io_y_sr = frontend_tlb_entries_barrier_5_io_y_sr;
    assign frontend_tlb__entries_barrier_5_io_y_hw = frontend_tlb_entries_barrier_5_io_y_hw;
    assign frontend_tlb__entries_barrier_5_io_y_hx = frontend_tlb_entries_barrier_5_io_y_hx;
    assign frontend_tlb__entries_barrier_5_io_y_hr = frontend_tlb_entries_barrier_5_io_y_hr;
     
  assign  frontend_tlb_io_resp_paddr ={ frontend_tlb_ppn , frontend_tlb_io_resp_gpa_offset }; 
  assign  frontend_tlb_io_resp_gpa ={ frontend_tlb_io_resp_gpa_page [19:0], frontend_tlb_io_resp_gpa_offset }; 
  assign  frontend_tlb_io_resp_pf_ld = frontend_tlb_pf_ld_array [6]; 
  assign  frontend_tlb_io_resp_pf_inst = frontend_tlb_pf_inst_array [6]; 
  assign  frontend_tlb_io_resp_ae_ld = frontend_tlb_ae_ld_array [6]; 
  assign  frontend_tlb_io_resp_ae_inst =~( frontend_tlb_px_array [6]); 
  assign  frontend_tlb_io_resp_ma_ld = frontend_tlb_misaligned ; 
  assign  frontend_tlb_io_resp_cacheable = frontend_tlb_c_array [6]; 
  assign  frontend_tlb_io_resp_prefetchable = frontend_tlb_prefetchable_array [6]; 
  assign  frontend_tlb_io_ptw_req_bits_valid =~ frontend_tlb_io_kill ; 
  assign  frontend_tlb_io_ptw_req_bits_bits_addr =20'h0; 
  assign  frontend_tlb_io_ptw_req_bits_bits_need_gpa =1'h0; 
  assign  frontend_tlb_io_ptw_req_bits_bits_vstage1 =1'h0; 
  assign  frontend_tlb_io_ptw_req_bits_bits_stage2 =1'h0;
    assign frontend_tlb_io_req_bits_vaddr = frontend_s1_pc;
    assign frontend__tlb_io_resp_paddr = frontend_tlb_io_resp_paddr;
    assign frontend__tlb_io_resp_gpa = frontend_tlb_io_resp_gpa;
    assign frontend__tlb_io_resp_pf_ld = frontend_tlb_io_resp_pf_ld;
    assign frontend__tlb_io_resp_pf_inst = frontend_tlb_io_resp_pf_inst;
    assign frontend__tlb_io_resp_ae_ld = frontend_tlb_io_resp_ae_ld;
    assign frontend__tlb_io_resp_ae_inst = frontend_tlb_io_resp_ae_inst;
    assign frontend__tlb_io_resp_ma_ld = frontend_tlb_io_resp_ma_ld;
    assign frontend__tlb_io_resp_cacheable = frontend_tlb_io_resp_cacheable;
    assign frontend__tlb_io_resp_prefetchable = frontend_tlb_io_resp_prefetchable;
    assign frontend_tlb_io_sfence_valid = frontend_io_cpu_sfence_valid;
    assign frontend_io_ptw_req_bits_valid = frontend_tlb_io_ptw_req_bits_valid;
    assign frontend_io_ptw_req_bits_bits_addr = frontend_tlb_io_ptw_req_bits_bits_addr;
    assign frontend_io_ptw_req_bits_bits_need_gpa = frontend_tlb_io_ptw_req_bits_bits_need_gpa;
    assign frontend_io_ptw_req_bits_bits_vstage1 = frontend_tlb_io_ptw_req_bits_bits_vstage1;
    assign frontend_io_ptw_req_bits_bits_stage2 = frontend_tlb_io_ptw_req_bits_bits_stage2;
    assign frontend_tlb_io_ptw_resp_bits_ae_ptw = frontend_io_ptw_resp_bits_ae_ptw;
    assign frontend_tlb_io_ptw_resp_bits_ae_final = frontend_io_ptw_resp_bits_ae_final;
    assign frontend_tlb_io_ptw_resp_bits_pf = frontend_io_ptw_resp_bits_pf;
    assign frontend_tlb_io_ptw_resp_bits_gf = frontend_io_ptw_resp_bits_gf;
    assign frontend_tlb_io_ptw_resp_bits_hr = frontend_io_ptw_resp_bits_hr;
    assign frontend_tlb_io_ptw_resp_bits_hw = frontend_io_ptw_resp_bits_hw;
    assign frontend_tlb_io_ptw_resp_bits_hx = frontend_io_ptw_resp_bits_hx;
    assign frontend_tlb_io_ptw_resp_bits_pte_ppn = frontend_io_ptw_resp_bits_pte_ppn;
    assign frontend_tlb_io_ptw_resp_bits_pte_d = frontend_io_ptw_resp_bits_pte_d;
    assign frontend_tlb_io_ptw_resp_bits_pte_a = frontend_io_ptw_resp_bits_pte_a;
    assign frontend_tlb_io_ptw_resp_bits_pte_g = frontend_io_ptw_resp_bits_pte_g;
    assign frontend_tlb_io_ptw_resp_bits_pte_u = frontend_io_ptw_resp_bits_pte_u;
    assign frontend_tlb_io_ptw_resp_bits_pte_x = frontend_io_ptw_resp_bits_pte_x;
    assign frontend_tlb_io_ptw_resp_bits_pte_w = frontend_io_ptw_resp_bits_pte_w;
    assign frontend_tlb_io_ptw_resp_bits_pte_r = frontend_io_ptw_resp_bits_pte_r;
    assign frontend_tlb_io_ptw_resp_bits_pte_v = frontend_io_ptw_resp_bits_pte_v;
    assign frontend_tlb_io_ptw_resp_bits_gpa_is_pte = frontend_io_ptw_resp_bits_gpa_is_pte;
    assign frontend_tlb_io_ptw_status_debug = frontend_io_ptw_status_debug;
    assign frontend_tlb_io_ptw_pmp_0_cfg_l = frontend_io_ptw_pmp_0_cfg_l;
    assign frontend_tlb_io_ptw_pmp_0_cfg_a = frontend_io_ptw_pmp_0_cfg_a;
    assign frontend_tlb_io_ptw_pmp_0_cfg_x = frontend_io_ptw_pmp_0_cfg_x;
    assign frontend_tlb_io_ptw_pmp_0_cfg_w = frontend_io_ptw_pmp_0_cfg_w;
    assign frontend_tlb_io_ptw_pmp_0_cfg_r = frontend_io_ptw_pmp_0_cfg_r;
    assign frontend_tlb_io_ptw_pmp_0_addr = frontend_io_ptw_pmp_0_addr;
    assign frontend_tlb_io_ptw_pmp_0_mask = frontend_io_ptw_pmp_0_mask;
    assign frontend_tlb_io_ptw_pmp_1_cfg_l = frontend_io_ptw_pmp_1_cfg_l;
    assign frontend_tlb_io_ptw_pmp_1_cfg_a = frontend_io_ptw_pmp_1_cfg_a;
    assign frontend_tlb_io_ptw_pmp_1_cfg_x = frontend_io_ptw_pmp_1_cfg_x;
    assign frontend_tlb_io_ptw_pmp_1_cfg_w = frontend_io_ptw_pmp_1_cfg_w;
    assign frontend_tlb_io_ptw_pmp_1_cfg_r = frontend_io_ptw_pmp_1_cfg_r;
    assign frontend_tlb_io_ptw_pmp_1_addr = frontend_io_ptw_pmp_1_addr;
    assign frontend_tlb_io_ptw_pmp_1_mask = frontend_io_ptw_pmp_1_mask;
    assign frontend_tlb_io_ptw_pmp_2_cfg_l = frontend_io_ptw_pmp_2_cfg_l;
    assign frontend_tlb_io_ptw_pmp_2_cfg_a = frontend_io_ptw_pmp_2_cfg_a;
    assign frontend_tlb_io_ptw_pmp_2_cfg_x = frontend_io_ptw_pmp_2_cfg_x;
    assign frontend_tlb_io_ptw_pmp_2_cfg_w = frontend_io_ptw_pmp_2_cfg_w;
    assign frontend_tlb_io_ptw_pmp_2_cfg_r = frontend_io_ptw_pmp_2_cfg_r;
    assign frontend_tlb_io_ptw_pmp_2_addr = frontend_io_ptw_pmp_2_addr;
    assign frontend_tlb_io_ptw_pmp_2_mask = frontend_io_ptw_pmp_2_mask;
    assign frontend_tlb_io_ptw_pmp_3_cfg_l = frontend_io_ptw_pmp_3_cfg_l;
    assign frontend_tlb_io_ptw_pmp_3_cfg_a = frontend_io_ptw_pmp_3_cfg_a;
    assign frontend_tlb_io_ptw_pmp_3_cfg_x = frontend_io_ptw_pmp_3_cfg_x;
    assign frontend_tlb_io_ptw_pmp_3_cfg_w = frontend_io_ptw_pmp_3_cfg_w;
    assign frontend_tlb_io_ptw_pmp_3_cfg_r = frontend_io_ptw_pmp_3_cfg_r;
    assign frontend_tlb_io_ptw_pmp_3_addr = frontend_io_ptw_pmp_3_addr;
    assign frontend_tlb_io_ptw_pmp_3_mask = frontend_io_ptw_pmp_3_mask;
    assign frontend_tlb_io_ptw_pmp_4_cfg_l = frontend_io_ptw_pmp_4_cfg_l;
    assign frontend_tlb_io_ptw_pmp_4_cfg_a = frontend_io_ptw_pmp_4_cfg_a;
    assign frontend_tlb_io_ptw_pmp_4_cfg_x = frontend_io_ptw_pmp_4_cfg_x;
    assign frontend_tlb_io_ptw_pmp_4_cfg_w = frontend_io_ptw_pmp_4_cfg_w;
    assign frontend_tlb_io_ptw_pmp_4_cfg_r = frontend_io_ptw_pmp_4_cfg_r;
    assign frontend_tlb_io_ptw_pmp_4_addr = frontend_io_ptw_pmp_4_addr;
    assign frontend_tlb_io_ptw_pmp_4_mask = frontend_io_ptw_pmp_4_mask;
    assign frontend_tlb_io_ptw_pmp_5_cfg_l = frontend_io_ptw_pmp_5_cfg_l;
    assign frontend_tlb_io_ptw_pmp_5_cfg_a = frontend_io_ptw_pmp_5_cfg_a;
    assign frontend_tlb_io_ptw_pmp_5_cfg_x = frontend_io_ptw_pmp_5_cfg_x;
    assign frontend_tlb_io_ptw_pmp_5_cfg_w = frontend_io_ptw_pmp_5_cfg_w;
    assign frontend_tlb_io_ptw_pmp_5_cfg_r = frontend_io_ptw_pmp_5_cfg_r;
    assign frontend_tlb_io_ptw_pmp_5_addr = frontend_io_ptw_pmp_5_addr;
    assign frontend_tlb_io_ptw_pmp_5_mask = frontend_io_ptw_pmp_5_mask;
    assign frontend_tlb_io_ptw_pmp_6_cfg_l = frontend_io_ptw_pmp_6_cfg_l;
    assign frontend_tlb_io_ptw_pmp_6_cfg_a = frontend_io_ptw_pmp_6_cfg_a;
    assign frontend_tlb_io_ptw_pmp_6_cfg_x = frontend_io_ptw_pmp_6_cfg_x;
    assign frontend_tlb_io_ptw_pmp_6_cfg_w = frontend_io_ptw_pmp_6_cfg_w;
    assign frontend_tlb_io_ptw_pmp_6_cfg_r = frontend_io_ptw_pmp_6_cfg_r;
    assign frontend_tlb_io_ptw_pmp_6_addr = frontend_io_ptw_pmp_6_addr;
    assign frontend_tlb_io_ptw_pmp_6_mask = frontend_io_ptw_pmp_6_mask;
    assign frontend_tlb_io_ptw_pmp_7_cfg_l = frontend_io_ptw_pmp_7_cfg_l;
    assign frontend_tlb_io_ptw_pmp_7_cfg_a = frontend_io_ptw_pmp_7_cfg_a;
    assign frontend_tlb_io_ptw_pmp_7_cfg_x = frontend_io_ptw_pmp_7_cfg_x;
    assign frontend_tlb_io_ptw_pmp_7_cfg_w = frontend_io_ptw_pmp_7_cfg_w;
    assign frontend_tlb_io_ptw_pmp_7_cfg_r = frontend_io_ptw_pmp_7_cfg_r;
    assign frontend_tlb_io_ptw_pmp_7_addr = frontend_io_ptw_pmp_7_addr;
    assign frontend_tlb_io_ptw_pmp_7_mask = frontend_io_ptw_pmp_7_mask;
    assign frontend_tlb_io_kill = ~frontend_s2_valid|frontend_s2_kill_speculative_tlb_refill;
     
  assign  frontend_io_cpu_gpa_valid = frontend_gpa_valid ; 
  assign  frontend_io_cpu_gpa_bits = frontend_gpa ;
    assign frontend_clock = clock;
    assign frontend_reset = reset;
    assign frontend_auto_icache_master_out_a_ready = widget_1_nodeIn_a_ready;
    assign widget_1_nodeIn_a_valid = frontend_auto_icache_master_out_a_valid;
    assign widget_1_nodeIn_a_bits_address = frontend_auto_icache_master_out_a_bits_address;
    assign widget_1_nodeIn_a_bits_user_amba_prot_readalloc = frontend_auto_icache_master_out_a_bits_user_amba_prot_readalloc;
    assign widget_1_nodeIn_a_bits_user_amba_prot_writealloc = frontend_auto_icache_master_out_a_bits_user_amba_prot_writealloc;
    assign frontend_auto_icache_master_out_d_valid = widget_1_nodeIn_d_valid;
    assign frontend_auto_icache_master_out_d_bits_opcode = widget_1_nodeIn_d_bits_opcode;
    assign frontend_auto_icache_master_out_d_bits_param = widget_1_nodeIn_d_bits_param;
    assign frontend_auto_icache_master_out_d_bits_size = widget_1_nodeIn_d_bits_size;
    assign frontend_auto_icache_master_out_d_bits_sink = widget_1_nodeIn_d_bits_sink;
    assign frontend_auto_icache_master_out_d_bits_denied = widget_1_nodeIn_d_bits_denied;
    assign frontend_auto_icache_master_out_d_bits_data = widget_1_nodeIn_d_bits_data;
    assign frontend_auto_icache_master_out_d_bits_corrupt = widget_1_nodeIn_d_bits_corrupt;
    assign frontend_io_cpu_might_request = _core_io_imem_might_request;
    assign frontend_io_cpu_req_valid = _core_io_imem_req_valid;
    assign frontend_io_cpu_req_bits_pc = _core_io_imem_req_bits_pc;
    assign frontend_io_cpu_req_bits_speculative = _core_io_imem_req_bits_speculative;
    assign frontend_io_cpu_sfence_valid = _core_io_imem_sfence_valid;
    assign frontend_io_cpu_resp_ready = _core_io_imem_resp_ready;
    assign _frontend_io_cpu_resp_valid = frontend_io_cpu_resp_valid;
    assign _frontend_io_cpu_resp_bits_btb_cfiType = frontend_io_cpu_resp_bits_btb_cfiType;
    assign _frontend_io_cpu_resp_bits_btb_taken = frontend_io_cpu_resp_bits_btb_taken;
    assign _frontend_io_cpu_resp_bits_btb_mask = frontend_io_cpu_resp_bits_btb_mask;
    assign _frontend_io_cpu_resp_bits_btb_bridx = frontend_io_cpu_resp_bits_btb_bridx;
    assign _frontend_io_cpu_resp_bits_btb_target = frontend_io_cpu_resp_bits_btb_target;
    assign _frontend_io_cpu_resp_bits_btb_entry = frontend_io_cpu_resp_bits_btb_entry;
    assign _frontend_io_cpu_resp_bits_btb_bht_history = frontend_io_cpu_resp_bits_btb_bht_history;
    assign _frontend_io_cpu_resp_bits_btb_bht_value = frontend_io_cpu_resp_bits_btb_bht_value;
    assign _frontend_io_cpu_resp_bits_pc = frontend_io_cpu_resp_bits_pc;
    assign _frontend_io_cpu_resp_bits_data = frontend_io_cpu_resp_bits_data;
    assign _frontend_io_cpu_resp_bits_mask = frontend_io_cpu_resp_bits_mask;
    assign _frontend_io_cpu_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst;
    assign _frontend_io_cpu_resp_bits_xcpt_gf_inst = frontend_io_cpu_resp_bits_xcpt_gf_inst;
    assign _frontend_io_cpu_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst;
    assign _frontend_io_cpu_resp_bits_replay = frontend_io_cpu_resp_bits_replay;
    assign _frontend_io_cpu_gpa_valid = frontend_io_cpu_gpa_valid;
    assign _frontend_io_cpu_gpa_bits = frontend_io_cpu_gpa_bits;
    assign frontend_io_cpu_btb_update_valid = _core_io_imem_btb_update_valid;
    assign frontend_io_cpu_bht_update_valid = _core_io_imem_bht_update_valid;
    assign frontend_io_cpu_flush_icache = _core_io_imem_flush_icache;
    assign frontend_io_cpu_progress = _core_io_imem_progress;
    assign _frontend_io_ptw_req_bits_valid = frontend_io_ptw_req_bits_valid;
    assign _frontend_io_ptw_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr;
    assign _frontend_io_ptw_req_bits_bits_need_gpa = frontend_io_ptw_req_bits_bits_need_gpa;
    assign _frontend_io_ptw_req_bits_bits_vstage1 = frontend_io_ptw_req_bits_bits_vstage1;
    assign _frontend_io_ptw_req_bits_bits_stage2 = frontend_io_ptw_req_bits_bits_stage2;
    assign frontend_io_ptw_resp_bits_ae_ptw = _ptw_io_requestor_1_resp_bits_ae_ptw;
    assign frontend_io_ptw_resp_bits_ae_final = _ptw_io_requestor_1_resp_bits_ae_final;
    assign frontend_io_ptw_resp_bits_pf = _ptw_io_requestor_1_resp_bits_pf;
    assign frontend_io_ptw_resp_bits_gf = _ptw_io_requestor_1_resp_bits_gf;
    assign frontend_io_ptw_resp_bits_hr = _ptw_io_requestor_1_resp_bits_hr;
    assign frontend_io_ptw_resp_bits_hw = _ptw_io_requestor_1_resp_bits_hw;
    assign frontend_io_ptw_resp_bits_hx = _ptw_io_requestor_1_resp_bits_hx;
    assign frontend_io_ptw_resp_bits_pte_ppn = _ptw_io_requestor_1_resp_bits_pte_ppn;
    assign frontend_io_ptw_resp_bits_pte_d = _ptw_io_requestor_1_resp_bits_pte_d;
    assign frontend_io_ptw_resp_bits_pte_a = _ptw_io_requestor_1_resp_bits_pte_a;
    assign frontend_io_ptw_resp_bits_pte_g = _ptw_io_requestor_1_resp_bits_pte_g;
    assign frontend_io_ptw_resp_bits_pte_u = _ptw_io_requestor_1_resp_bits_pte_u;
    assign frontend_io_ptw_resp_bits_pte_x = _ptw_io_requestor_1_resp_bits_pte_x;
    assign frontend_io_ptw_resp_bits_pte_w = _ptw_io_requestor_1_resp_bits_pte_w;
    assign frontend_io_ptw_resp_bits_pte_r = _ptw_io_requestor_1_resp_bits_pte_r;
    assign frontend_io_ptw_resp_bits_pte_v = _ptw_io_requestor_1_resp_bits_pte_v;
    assign frontend_io_ptw_resp_bits_gpa_is_pte = _ptw_io_requestor_1_resp_bits_gpa_is_pte;
    assign frontend_io_ptw_status_debug = _ptw_io_requestor_1_status_debug;
    assign frontend_io_ptw_pmp_0_cfg_l = _ptw_io_requestor_1_pmp_0_cfg_l;
    assign frontend_io_ptw_pmp_0_cfg_a = _ptw_io_requestor_1_pmp_0_cfg_a;
    assign frontend_io_ptw_pmp_0_cfg_x = _ptw_io_requestor_1_pmp_0_cfg_x;
    assign frontend_io_ptw_pmp_0_cfg_w = _ptw_io_requestor_1_pmp_0_cfg_w;
    assign frontend_io_ptw_pmp_0_cfg_r = _ptw_io_requestor_1_pmp_0_cfg_r;
    assign frontend_io_ptw_pmp_0_addr = _ptw_io_requestor_1_pmp_0_addr;
    assign frontend_io_ptw_pmp_0_mask = _ptw_io_requestor_1_pmp_0_mask;
    assign frontend_io_ptw_pmp_1_cfg_l = _ptw_io_requestor_1_pmp_1_cfg_l;
    assign frontend_io_ptw_pmp_1_cfg_a = _ptw_io_requestor_1_pmp_1_cfg_a;
    assign frontend_io_ptw_pmp_1_cfg_x = _ptw_io_requestor_1_pmp_1_cfg_x;
    assign frontend_io_ptw_pmp_1_cfg_w = _ptw_io_requestor_1_pmp_1_cfg_w;
    assign frontend_io_ptw_pmp_1_cfg_r = _ptw_io_requestor_1_pmp_1_cfg_r;
    assign frontend_io_ptw_pmp_1_addr = _ptw_io_requestor_1_pmp_1_addr;
    assign frontend_io_ptw_pmp_1_mask = _ptw_io_requestor_1_pmp_1_mask;
    assign frontend_io_ptw_pmp_2_cfg_l = _ptw_io_requestor_1_pmp_2_cfg_l;
    assign frontend_io_ptw_pmp_2_cfg_a = _ptw_io_requestor_1_pmp_2_cfg_a;
    assign frontend_io_ptw_pmp_2_cfg_x = _ptw_io_requestor_1_pmp_2_cfg_x;
    assign frontend_io_ptw_pmp_2_cfg_w = _ptw_io_requestor_1_pmp_2_cfg_w;
    assign frontend_io_ptw_pmp_2_cfg_r = _ptw_io_requestor_1_pmp_2_cfg_r;
    assign frontend_io_ptw_pmp_2_addr = _ptw_io_requestor_1_pmp_2_addr;
    assign frontend_io_ptw_pmp_2_mask = _ptw_io_requestor_1_pmp_2_mask;
    assign frontend_io_ptw_pmp_3_cfg_l = _ptw_io_requestor_1_pmp_3_cfg_l;
    assign frontend_io_ptw_pmp_3_cfg_a = _ptw_io_requestor_1_pmp_3_cfg_a;
    assign frontend_io_ptw_pmp_3_cfg_x = _ptw_io_requestor_1_pmp_3_cfg_x;
    assign frontend_io_ptw_pmp_3_cfg_w = _ptw_io_requestor_1_pmp_3_cfg_w;
    assign frontend_io_ptw_pmp_3_cfg_r = _ptw_io_requestor_1_pmp_3_cfg_r;
    assign frontend_io_ptw_pmp_3_addr = _ptw_io_requestor_1_pmp_3_addr;
    assign frontend_io_ptw_pmp_3_mask = _ptw_io_requestor_1_pmp_3_mask;
    assign frontend_io_ptw_pmp_4_cfg_l = _ptw_io_requestor_1_pmp_4_cfg_l;
    assign frontend_io_ptw_pmp_4_cfg_a = _ptw_io_requestor_1_pmp_4_cfg_a;
    assign frontend_io_ptw_pmp_4_cfg_x = _ptw_io_requestor_1_pmp_4_cfg_x;
    assign frontend_io_ptw_pmp_4_cfg_w = _ptw_io_requestor_1_pmp_4_cfg_w;
    assign frontend_io_ptw_pmp_4_cfg_r = _ptw_io_requestor_1_pmp_4_cfg_r;
    assign frontend_io_ptw_pmp_4_addr = _ptw_io_requestor_1_pmp_4_addr;
    assign frontend_io_ptw_pmp_4_mask = _ptw_io_requestor_1_pmp_4_mask;
    assign frontend_io_ptw_pmp_5_cfg_l = _ptw_io_requestor_1_pmp_5_cfg_l;
    assign frontend_io_ptw_pmp_5_cfg_a = _ptw_io_requestor_1_pmp_5_cfg_a;
    assign frontend_io_ptw_pmp_5_cfg_x = _ptw_io_requestor_1_pmp_5_cfg_x;
    assign frontend_io_ptw_pmp_5_cfg_w = _ptw_io_requestor_1_pmp_5_cfg_w;
    assign frontend_io_ptw_pmp_5_cfg_r = _ptw_io_requestor_1_pmp_5_cfg_r;
    assign frontend_io_ptw_pmp_5_addr = _ptw_io_requestor_1_pmp_5_addr;
    assign frontend_io_ptw_pmp_5_mask = _ptw_io_requestor_1_pmp_5_mask;
    assign frontend_io_ptw_pmp_6_cfg_l = _ptw_io_requestor_1_pmp_6_cfg_l;
    assign frontend_io_ptw_pmp_6_cfg_a = _ptw_io_requestor_1_pmp_6_cfg_a;
    assign frontend_io_ptw_pmp_6_cfg_x = _ptw_io_requestor_1_pmp_6_cfg_x;
    assign frontend_io_ptw_pmp_6_cfg_w = _ptw_io_requestor_1_pmp_6_cfg_w;
    assign frontend_io_ptw_pmp_6_cfg_r = _ptw_io_requestor_1_pmp_6_cfg_r;
    assign frontend_io_ptw_pmp_6_addr = _ptw_io_requestor_1_pmp_6_addr;
    assign frontend_io_ptw_pmp_6_mask = _ptw_io_requestor_1_pmp_6_mask;
    assign frontend_io_ptw_pmp_7_cfg_l = _ptw_io_requestor_1_pmp_7_cfg_l;
    assign frontend_io_ptw_pmp_7_cfg_a = _ptw_io_requestor_1_pmp_7_cfg_a;
    assign frontend_io_ptw_pmp_7_cfg_x = _ptw_io_requestor_1_pmp_7_cfg_x;
    assign frontend_io_ptw_pmp_7_cfg_w = _ptw_io_requestor_1_pmp_7_cfg_w;
    assign frontend_io_ptw_pmp_7_cfg_r = _ptw_io_requestor_1_pmp_7_cfg_r;
    assign frontend_io_ptw_pmp_7_addr = _ptw_io_requestor_1_pmp_7_addr;
    assign frontend_io_ptw_pmp_7_mask = _ptw_io_requestor_1_pmp_7_mask;
    assign frontend_io_ptw_customCSRs_csrs_0_value = _ptw_io_requestor_1_customCSRs_csrs_0_value;
    
  wire dtim_adapter_clock;
    wire dtim_adapter_reset;
    wire dtim_adapter_auto_in_a_ready;
    wire dtim_adapter_auto_in_a_valid;
    wire[2:0] dtim_adapter_auto_in_a_bits_opcode;
    wire[2:0] dtim_adapter_auto_in_a_bits_param;
    wire[1:0] dtim_adapter_auto_in_a_bits_size;
    wire[10:0] dtim_adapter_auto_in_a_bits_source;
    wire[31:0] dtim_adapter_auto_in_a_bits_address;
    wire[3:0] dtim_adapter_auto_in_a_bits_mask;
    wire[31:0] dtim_adapter_auto_in_a_bits_data;
    wire dtim_adapter_auto_in_a_bits_corrupt;
    wire dtim_adapter_auto_in_d_ready;
    wire dtim_adapter_auto_in_d_valid;
    wire[2:0] dtim_adapter_auto_in_d_bits_opcode;
    wire[1:0] dtim_adapter_auto_in_d_bits_size;
    wire[10:0] dtim_adapter_auto_in_d_bits_source;
    wire[31:0] dtim_adapter_auto_in_d_bits_data;
    wire dtim_adapter_io_dmem_req_ready;
    wire dtim_adapter_io_dmem_req_valid;
    wire[31:0] dtim_adapter_io_dmem_req_bits_addr;
    wire[4:0] dtim_adapter_io_dmem_req_bits_cmd;
    wire[1:0] dtim_adapter_io_dmem_req_bits_size;
    wire dtim_adapter_io_dmem_s1_kill;
    wire[31:0] dtim_adapter_io_dmem_s1_data_data;
    wire[3:0] dtim_adapter_io_dmem_s1_data_mask;
    wire dtim_adapter_io_dmem_s2_nack;
    wire dtim_adapter_io_dmem_resp_valid;
    wire[31:0] dtim_adapter_io_dmem_resp_bits_data_raw;

    wire dtim_adapter_nodeIn_a_valid = dtim_adapter_auto_in_a_valid ; 
    wire[2:0] dtim_adapter_nodeIn_a_bits_opcode = dtim_adapter_auto_in_a_bits_opcode ; 
    wire[2:0] dtim_adapter_nodeIn_a_bits_param = dtim_adapter_auto_in_a_bits_param ; 
    wire[1:0] dtim_adapter_nodeIn_a_bits_size = dtim_adapter_auto_in_a_bits_size ; 
    wire[10:0] dtim_adapter_nodeIn_a_bits_source = dtim_adapter_auto_in_a_bits_source ; 
    wire[31:0] dtim_adapter_nodeIn_a_bits_address = dtim_adapter_auto_in_a_bits_address ; 
    wire[3:0] dtim_adapter_nodeIn_a_bits_mask = dtim_adapter_auto_in_a_bits_mask ; 
    wire[31:0] dtim_adapter_nodeIn_a_bits_data = dtim_adapter_auto_in_a_bits_data ; 
    wire dtim_adapter_nodeIn_a_bits_corrupt = dtim_adapter_auto_in_a_bits_corrupt ; 
    wire dtim_adapter_nodeIn_d_ready = dtim_adapter_auto_in_d_ready ; 
    wire[1:0] dtim_adapter_nodeIn_d_bits_param =2'h0; 
    wire[1:0] dtim_adapter_io_dmem_req_bits_req_dprv =2'h0; 
    wire[1:0] dtim_adapter_nodeIn_d_bits_d_param =2'h0; 
    wire[1:0] dtim_adapter_nodeIn_d_bits_d_1_param =2'h0; 
    wire dtim_adapter_io_dmem_req_bits_req_phys =1'h1; 
    wire dtim_adapter_io_dmem_req_bits_req_no_xcpt =1'h1; 
    wire[6:0] dtim_adapter_io_dmem_req_bits_req_tag =7'h0; 
    wire[3:0] dtim_adapter_io_dmem_req_bits_req_mask =4'h0; 
    wire[31:0] dtim_adapter_io_dmem_req_bits_req_data =32'h0; 
    wire[31:0] dtim_adapter_nodeIn_d_bits_d_data =32'h0; 
    wire[31:0] dtim_adapter_nodeIn_d_bits_d_1_data =32'h0; 
    wire[2:0] dtim_adapter_nodeIn_d_bits_d_opcode =3'h0; 
    wire[2:0] dtim_adapter_nodeIn_d_bits_d_1_opcode =3'h1; 
    wire dtim_adapter_nodeIn_d_bits_sink =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_denied =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_corrupt =1'h0; 
    wire dtim_adapter_io_dmem_req_bits_req_signed =1'h0; 
    wire dtim_adapter_io_dmem_req_bits_req_dv =1'h0; 
    wire dtim_adapter_io_dmem_req_bits_req_no_alloc =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_d_sink =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_d_denied =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_d_corrupt =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_d_1_sink =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_d_1_denied =1'h0; 
    wire dtim_adapter_nodeIn_d_bits_d_1_corrupt =1'h0; reg[2:0] dtim_adapter_state ; 
    wire dtim_adapter__io_dmem_req_bits_T_2 = dtim_adapter_state ==3'h4; reg[2:0] dtim_adapter_acq_opcode ; reg[2:0] dtim_adapter_acq_param ; reg[1:0] dtim_adapter_acq_size ; 
    wire[1:0] dtim_adapter_nodeIn_d_bits_d_size = dtim_adapter_acq_size ; 
    wire[1:0] dtim_adapter_nodeIn_d_bits_d_1_size = dtim_adapter_acq_size ; reg[10:0] dtim_adapter_acq_source ; 
    wire[10:0] dtim_adapter_nodeIn_d_bits_d_source = dtim_adapter_acq_source ; 
    wire[10:0] dtim_adapter_nodeIn_d_bits_d_1_source = dtim_adapter_acq_source ; reg[31:0] dtim_adapter_acq_address ; reg[3:0] dtim_adapter_acq_mask ; reg[31:0] dtim_adapter_acq_data ; 
    reg dtim_adapter_acq_corrupt ; 
    wire dtim_adapter__ready_T = dtim_adapter_state ==3'h0; 
    wire dtim_adapter__nodeIn_d_bits_data_T = dtim_adapter_state ==3'h2; 
    wire dtim_adapter_ready_likely = dtim_adapter__ready_T | dtim_adapter__nodeIn_d_bits_data_T ; 
    wire dtim_adapter_ready = dtim_adapter__ready_T | dtim_adapter__nodeIn_d_bits_data_T & dtim_adapter_io_dmem_resp_valid & dtim_adapter_nodeIn_d_ready ; 
    wire dtim_adapter__io_dmem_req_bits_T = dtim_adapter_state ==3'h3; 
    wire dtim_adapter_dmem_req_valid = dtim_adapter_nodeIn_a_valid & dtim_adapter_ready | dtim_adapter__io_dmem_req_bits_T ; 
    wire dtim_adapter_dmem_req_valid_likely = dtim_adapter_nodeIn_a_valid & dtim_adapter_ready_likely | dtim_adapter__io_dmem_req_bits_T ; 
    wire dtim_adapter_nodeIn_a_ready = dtim_adapter_io_dmem_req_ready & dtim_adapter_ready ; 
    wire[2:0] dtim_adapter__io_dmem_req_bits_T_1_opcode = dtim_adapter__io_dmem_req_bits_T  ?  dtim_adapter_acq_opcode : dtim_adapter_nodeIn_a_bits_opcode ; 
    wire[2:0] dtim_adapter__io_dmem_req_bits_T_1_param = dtim_adapter__io_dmem_req_bits_T  ?  dtim_adapter_acq_param : dtim_adapter_nodeIn_a_bits_param ; 
    wire[1:0] dtim_adapter__io_dmem_req_bits_T_1_size = dtim_adapter__io_dmem_req_bits_T  ?  dtim_adapter_acq_size : dtim_adapter_nodeIn_a_bits_size ; 
    wire[1:0] dtim_adapter_io_dmem_req_bits_req_size ; 
  assign  dtim_adapter_io_dmem_req_bits_req_size = dtim_adapter__io_dmem_req_bits_T_1_size ; 
    wire[1:0] dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_size ; 
  assign  dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_size = dtim_adapter__io_dmem_req_bits_T_1_size ; 
    wire[31:0] dtim_adapter_io_dmem_req_bits_req_addr = dtim_adapter__io_dmem_req_bits_T  ?  dtim_adapter_acq_address : dtim_adapter_nodeIn_a_bits_address ; reg[3:0] dtim_adapter_casez_tmp ; 
  always @(*)
         begin 
             casez ( dtim_adapter__io_dmem_req_bits_T_1_param )
              3 'b000: 
                  dtim_adapter_casez_tmp  =4'hC;
              3 'b001: 
                  dtim_adapter_casez_tmp  =4'hD;
              3 'b010: 
                  dtim_adapter_casez_tmp  =4'hE;
              3 'b011: 
                  dtim_adapter_casez_tmp  =4'hF;
              3 'b100: 
                  dtim_adapter_casez_tmp  =4'h8;
              3 'b101: 
                  dtim_adapter_casez_tmp  =4'h0;
              3 'b110: 
                  dtim_adapter_casez_tmp  =4'h0;
              default : 
                  dtim_adapter_casez_tmp  =4'h0;endcase
         end
    wire dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_upper = dtim_adapter_io_dmem_req_bits_req_addr [0]|(| dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_size ); 
    wire dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_lower =~( dtim_adapter_io_dmem_req_bits_req_addr [0]); 
    wire[1:0] dtim_adapter__io_dmem_req_bits_mask_full_desired_mask_T ={ dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_upper , dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_lower }; 
    wire[1:0] dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_upper_1 =( dtim_adapter_io_dmem_req_bits_req_addr [1] ?  dtim_adapter__io_dmem_req_bits_mask_full_desired_mask_T :2'h0)|{2{ dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_size [1]}}; 
    wire[1:0] dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_lower_1 = dtim_adapter_io_dmem_req_bits_req_addr [1] ? 2'h0: dtim_adapter__io_dmem_req_bits_mask_full_desired_mask_T ; 
    wire[3:0] dtim_adapter_io_dmem_req_bits_mask_full_desired_mask ={ dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_upper_1 , dtim_adapter_io_dmem_req_bits_mask_full_desired_mask_lower_1 }; 
    wire dtim_adapter_io_dmem_req_bits_mask_full =&(( dtim_adapter__io_dmem_req_bits_T  ?  dtim_adapter_acq_mask : dtim_adapter_nodeIn_a_bits_mask )|~ dtim_adapter_io_dmem_req_bits_mask_full_desired_mask ); 
    wire[4:0] dtim_adapter_io_dmem_req_bits_req_cmd = dtim_adapter__io_dmem_req_bits_T_2 | dtim_adapter__io_dmem_req_bits_T_1_opcode ==3'h1& dtim_adapter_io_dmem_req_bits_mask_full  ? 5'h1: dtim_adapter__io_dmem_req_bits_T_1_opcode ==3'h4 ? 5'h0: dtim_adapter__io_dmem_req_bits_T_1_opcode ==3'h3 ? {1'h0, dtim_adapter__io_dmem_req_bits_T_1_param ==3'h3 ? 4'h4: dtim_adapter__io_dmem_req_bits_T_1_param ==3'h2 ? 4'hB: dtim_adapter__io_dmem_req_bits_T_1_param ==3'h1 ? 4'hA: dtim_adapter__io_dmem_req_bits_T_1_param ==3'h0 ? 4'h9:4'h0}: dtim_adapter__io_dmem_req_bits_T_1_opcode ==3'h2 ? {1'h0, dtim_adapter_casez_tmp }: dtim_adapter__io_dmem_req_bits_T_1_opcode ==3'h1 ? 5'h11:{4'h0, dtim_adapter__io_dmem_req_bits_T_1_opcode ==3'h0}; 
    wire dtim_adapter_nodeIn_d_valid = dtim_adapter_io_dmem_resp_valid | dtim_adapter_state ==3'h5; 
    wire dtim_adapter__nodeIn_d_bits_T_2 = dtim_adapter_acq_opcode ==3'h0| dtim_adapter_acq_opcode ==3'h1; 
    wire[2:0] dtim_adapter_nodeIn_d_bits_opcode ={2'h0,~ dtim_adapter__nodeIn_d_bits_T_2 }; 
    wire[1:0] dtim_adapter_nodeIn_d_bits_size = dtim_adapter__nodeIn_d_bits_T_2  ?  dtim_adapter_nodeIn_d_bits_d_size : dtim_adapter_nodeIn_d_bits_d_1_size ; 
    wire[10:0] dtim_adapter_nodeIn_d_bits_source = dtim_adapter__nodeIn_d_bits_T_2  ?  dtim_adapter_nodeIn_d_bits_d_source : dtim_adapter_nodeIn_d_bits_d_1_source ; reg[31:0] dtim_adapter_nodeIn_d_bits_data_r ; 
    wire[31:0] dtim_adapter_nodeIn_d_bits_data = dtim_adapter__nodeIn_d_bits_data_T  ?  dtim_adapter_io_dmem_resp_bits_data_raw : dtim_adapter_nodeIn_d_bits_data_r ; 
  always @( posedge  dtim_adapter_clock )
         begin 
             if ( dtim_adapter_reset ) 
                 dtim_adapter_state  <=3'h4;
              else 
                 if ( dtim_adapter_dmem_req_valid & dtim_adapter_io_dmem_req_ready ) 
                     dtim_adapter_state  <=3'h1;
                  else 
                     if ( dtim_adapter_io_dmem_s2_nack ) 
                         dtim_adapter_state  <=3'h3;
                      else 
                         if ( dtim_adapter_nodeIn_d_ready & dtim_adapter_nodeIn_d_valid ) 
                             dtim_adapter_state  <=3'h0;
                          else 
                             if ( dtim_adapter_io_dmem_resp_valid ) 
                                 dtim_adapter_state  <=3'h5;
                              else 
                                 if ( dtim_adapter__io_dmem_req_bits_T_2 & dtim_adapter_nodeIn_a_valid ) 
                                     dtim_adapter_state  <=3'h0;
                                  else 
                                     if ( dtim_adapter_state ==3'h1) 
                                         dtim_adapter_state  <=3'h2;
             if ( dtim_adapter_nodeIn_a_ready & dtim_adapter_nodeIn_a_valid )
                 begin  
                     dtim_adapter_acq_opcode  <= dtim_adapter_nodeIn_a_bits_opcode ; 
                     dtim_adapter_acq_param  <= dtim_adapter_nodeIn_a_bits_param ; 
                     dtim_adapter_acq_size  <= dtim_adapter_nodeIn_a_bits_size ; 
                     dtim_adapter_acq_source  <= dtim_adapter_nodeIn_a_bits_source ; 
                     dtim_adapter_acq_address  <= dtim_adapter_nodeIn_a_bits_address ; 
                     dtim_adapter_acq_mask  <= dtim_adapter_nodeIn_a_bits_mask ; 
                     dtim_adapter_acq_data  <= dtim_adapter_nodeIn_a_bits_data ; 
                     dtim_adapter_acq_corrupt  <= dtim_adapter_nodeIn_a_bits_corrupt ;
                 end 
             if ( dtim_adapter__nodeIn_d_bits_data_T ) 
                 dtim_adapter_nodeIn_d_bits_data_r  <= dtim_adapter_io_dmem_resp_bits_data_raw ;
         end
  assign  dtim_adapter_auto_in_a_ready = dtim_adapter_nodeIn_a_ready ; 
  assign  dtim_adapter_auto_in_d_valid = dtim_adapter_nodeIn_d_valid ; 
  assign  dtim_adapter_auto_in_d_bits_opcode = dtim_adapter_nodeIn_d_bits_opcode ; 
  assign  dtim_adapter_auto_in_d_bits_size = dtim_adapter_nodeIn_d_bits_size ; 
  assign  dtim_adapter_auto_in_d_bits_source = dtim_adapter_nodeIn_d_bits_source ; 
  assign  dtim_adapter_auto_in_d_bits_data = dtim_adapter_nodeIn_d_bits_data ; 
  assign  dtim_adapter_io_dmem_req_valid = dtim_adapter_dmem_req_valid_likely ; 
  assign  dtim_adapter_io_dmem_req_bits_addr = dtim_adapter_io_dmem_req_bits_req_addr ; 
  assign  dtim_adapter_io_dmem_req_bits_cmd = dtim_adapter_io_dmem_req_bits_req_cmd ; 
  assign  dtim_adapter_io_dmem_req_bits_size = dtim_adapter_io_dmem_req_bits_req_size ; 
  assign  dtim_adapter_io_dmem_s1_kill = dtim_adapter_state !=3'h1; 
  assign  dtim_adapter_io_dmem_s1_data_data = dtim_adapter_acq_data ; 
  assign  dtim_adapter_io_dmem_s1_data_mask = dtim_adapter_acq_mask ;
    assign dtim_adapter_clock = clock;
    assign dtim_adapter_reset = reset;
    assign _dtim_adapter_auto_in_a_ready = dtim_adapter_auto_in_a_ready;
    assign dtim_adapter_auto_in_a_valid = _fragmenter_1_auto_out_a_valid;
    assign dtim_adapter_auto_in_a_bits_opcode = _fragmenter_1_auto_out_a_bits_opcode;
    assign dtim_adapter_auto_in_a_bits_param = _fragmenter_1_auto_out_a_bits_param;
    assign dtim_adapter_auto_in_a_bits_size = _fragmenter_1_auto_out_a_bits_size;
    assign dtim_adapter_auto_in_a_bits_source = _fragmenter_1_auto_out_a_bits_source;
    assign dtim_adapter_auto_in_a_bits_address = _fragmenter_1_auto_out_a_bits_address;
    assign dtim_adapter_auto_in_a_bits_mask = _fragmenter_1_auto_out_a_bits_mask;
    assign dtim_adapter_auto_in_a_bits_data = _fragmenter_1_auto_out_a_bits_data;
    assign dtim_adapter_auto_in_a_bits_corrupt = _fragmenter_1_auto_out_a_bits_corrupt;
    assign dtim_adapter_auto_in_d_ready = _fragmenter_1_auto_out_d_ready;
    assign _dtim_adapter_auto_in_d_valid = dtim_adapter_auto_in_d_valid;
    assign _dtim_adapter_auto_in_d_bits_opcode = dtim_adapter_auto_in_d_bits_opcode;
    assign _dtim_adapter_auto_in_d_bits_size = dtim_adapter_auto_in_d_bits_size;
    assign _dtim_adapter_auto_in_d_bits_source = dtim_adapter_auto_in_d_bits_source;
    assign _dtim_adapter_auto_in_d_bits_data = dtim_adapter_auto_in_d_bits_data;
    assign dtim_adapter_io_dmem_req_ready = _dcacheArb_io_requestor_1_req_ready;
    assign _dtim_adapter_io_dmem_req_valid = dtim_adapter_io_dmem_req_valid;
    assign _dtim_adapter_io_dmem_req_bits_addr = dtim_adapter_io_dmem_req_bits_addr;
    assign _dtim_adapter_io_dmem_req_bits_cmd = dtim_adapter_io_dmem_req_bits_cmd;
    assign _dtim_adapter_io_dmem_req_bits_size = dtim_adapter_io_dmem_req_bits_size;
    assign _dtim_adapter_io_dmem_s1_kill = dtim_adapter_io_dmem_s1_kill;
    assign _dtim_adapter_io_dmem_s1_data_data = dtim_adapter_io_dmem_s1_data_data;
    assign _dtim_adapter_io_dmem_s1_data_mask = dtim_adapter_io_dmem_s1_data_mask;
    assign dtim_adapter_io_dmem_s2_nack = _dcacheArb_io_requestor_1_s2_nack;
    assign dtim_adapter_io_dmem_resp_valid = _dcacheArb_io_requestor_1_resp_valid;
    assign dtim_adapter_io_dmem_resp_bits_data_raw = _dcacheArb_io_requestor_1_resp_bits_data_raw;
    
  wire fragmenter_1_clock;
    wire fragmenter_1_reset;
    wire fragmenter_1_auto_in_a_ready;
    wire fragmenter_1_auto_in_a_valid;
    wire[2:0] fragmenter_1_auto_in_a_bits_opcode;
    wire[2:0] fragmenter_1_auto_in_a_bits_param;
    wire[2:0] fragmenter_1_auto_in_a_bits_size;
    wire[4:0] fragmenter_1_auto_in_a_bits_source;
    wire[31:0] fragmenter_1_auto_in_a_bits_address;
    wire[3:0] fragmenter_1_auto_in_a_bits_mask;
    wire[31:0] fragmenter_1_auto_in_a_bits_data;
    wire fragmenter_1_auto_in_a_bits_corrupt;
    wire fragmenter_1_auto_in_d_ready;
    wire fragmenter_1_auto_in_d_valid;
    wire[2:0] fragmenter_1_auto_in_d_bits_opcode;
    wire[2:0] fragmenter_1_auto_in_d_bits_size;
    wire[4:0] fragmenter_1_auto_in_d_bits_source;
    wire[31:0] fragmenter_1_auto_in_d_bits_data;
    wire fragmenter_1_auto_out_a_ready;
    wire fragmenter_1_auto_out_a_valid;
    wire[2:0] fragmenter_1_auto_out_a_bits_opcode;
    wire[2:0] fragmenter_1_auto_out_a_bits_param;
    wire[1:0] fragmenter_1_auto_out_a_bits_size;
    wire[10:0] fragmenter_1_auto_out_a_bits_source;
    wire[31:0] fragmenter_1_auto_out_a_bits_address;
    wire[3:0] fragmenter_1_auto_out_a_bits_mask;
    wire[31:0] fragmenter_1_auto_out_a_bits_data;
    wire fragmenter_1_auto_out_a_bits_corrupt;
    wire fragmenter_1_auto_out_d_ready;
    wire fragmenter_1_auto_out_d_valid;
    wire[2:0] fragmenter_1_auto_out_d_bits_opcode;
    wire[1:0] fragmenter_1_auto_out_d_bits_size;
    wire[10:0] fragmenter_1_auto_out_d_bits_source;
    wire[31:0] fragmenter_1_auto_out_d_bits_data;

    wire fragmenter_1_nodeOut_a_bits_corrupt ; 
    wire[2:0] fragmenter_1_nodeOut_a_bits_param ; 
    wire fragmenter_1_nodeIn_a_ready ; 
    wire fragmenter_1__repeater_io_full ; 
    wire[2:0] fragmenter_1__repeater_io_deq_bits_opcode ; 
    wire[2:0] fragmenter_1__repeater_io_deq_bits_size ; 
    wire[4:0] fragmenter_1__repeater_io_deq_bits_source ; 
    wire[31:0] fragmenter_1__repeater_io_deq_bits_address ; 
    wire[3:0] fragmenter_1__repeater_io_deq_bits_mask ; 
    wire fragmenter_1_nodeIn_a_valid = fragmenter_1_auto_in_a_valid ; 
    wire[2:0] fragmenter_1_nodeIn_a_bits_opcode = fragmenter_1_auto_in_a_bits_opcode ; 
    wire[2:0] fragmenter_1_nodeIn_a_bits_param = fragmenter_1_auto_in_a_bits_param ; 
    wire[2:0] fragmenter_1_nodeIn_a_bits_size = fragmenter_1_auto_in_a_bits_size ; 
    wire[4:0] fragmenter_1_nodeIn_a_bits_source = fragmenter_1_auto_in_a_bits_source ; 
    wire[31:0] fragmenter_1_nodeIn_a_bits_address = fragmenter_1_auto_in_a_bits_address ; 
    wire[3:0] fragmenter_1_nodeIn_a_bits_mask = fragmenter_1_auto_in_a_bits_mask ; 
    wire[31:0] fragmenter_1_nodeIn_a_bits_data = fragmenter_1_auto_in_a_bits_data ; 
    wire fragmenter_1_nodeIn_a_bits_corrupt = fragmenter_1_auto_in_a_bits_corrupt ; 
    wire fragmenter_1_nodeIn_d_ready = fragmenter_1_auto_in_d_ready ; 
    wire fragmenter_1_nodeOut_a_ready = fragmenter_1_auto_out_a_ready ; 
    wire fragmenter_1_nodeOut_d_valid = fragmenter_1_auto_out_d_valid ; 
    wire[2:0] fragmenter_1_nodeOut_d_bits_opcode = fragmenter_1_auto_out_d_bits_opcode ; 
    wire[1:0] fragmenter_1_nodeOut_d_bits_size = fragmenter_1_auto_out_d_bits_size ; 
    wire[10:0] fragmenter_1_nodeOut_d_bits_source = fragmenter_1_auto_out_d_bits_source ; 
    wire[31:0] fragmenter_1_nodeOut_d_bits_data = fragmenter_1_auto_out_d_bits_data ; 
    wire[1:0] fragmenter_1_nodeIn_d_bits_param =2'h0; 
    wire[1:0] fragmenter_1_nodeOut_d_bits_param =2'h0; 
    wire fragmenter_1_nodeIn_d_bits_sink =1'h0; 
    wire fragmenter_1_nodeIn_d_bits_denied =1'h0; 
    wire fragmenter_1_nodeIn_d_bits_corrupt =1'h0; 
    wire fragmenter_1_nodeOut_d_bits_sink =1'h0; 
    wire fragmenter_1_nodeOut_d_bits_denied =1'h0; 
    wire fragmenter_1_nodeOut_d_bits_corrupt =1'h0; 
    wire fragmenter_1_acknum_size =1'h0; 
    wire fragmenter_1_find_0 =1'h1; 
    wire[1:0] fragmenter_1_limit =2'h2; 
    wire[31:0] fragmenter_1_nodeOut_a_bits_data = fragmenter_1_nodeIn_a_bits_data ; 
    wire[2:0] fragmenter_1_nodeIn_d_bits_opcode = fragmenter_1_nodeOut_d_bits_opcode ; 
    wire[1:0] fragmenter_1_dsizeOH_shiftAmount = fragmenter_1_nodeOut_d_bits_size ; 
    wire[31:0] fragmenter_1_nodeIn_d_bits_data = fragmenter_1_nodeOut_d_bits_data ; reg[3:0] fragmenter_1_acknum ; reg[2:0] fragmenter_1_dOrig ; 
    reg fragmenter_1_dToggle ; 
    wire[3:0] fragmenter_1_dFragnum = fragmenter_1_nodeOut_d_bits_source [3:0]; 
    wire[3:0] fragmenter_1_acknum_fragment = fragmenter_1_dFragnum ; 
    wire fragmenter_1_dFirst = fragmenter_1_acknum ==4'h0; 
    wire fragmenter_1_dLast = fragmenter_1_dFragnum ==4'h0; 
    wire[3:0] fragmenter_1__dsizeOH_T =4'h1<< fragmenter_1_dsizeOH_shiftAmount ; 
    wire[2:0] fragmenter_1_dsizeOH = fragmenter_1__dsizeOH_T [2:0]; 
    wire[4:0] fragmenter_1__dsizeOH1_T_1 =5'h3<< fragmenter_1_nodeOut_d_bits_size ; 
    wire[1:0] fragmenter_1_dsizeOH1 =~( fragmenter_1__dsizeOH1_T_1 [1:0]); 
    wire fragmenter_1_dHasData = fragmenter_1_nodeOut_d_bits_opcode [0]; 
    wire[3:0] fragmenter_1_dFirst_acknum = fragmenter_1_acknum_fragment ; 
    wire fragmenter_1_ack_decrement = fragmenter_1_dHasData | fragmenter_1_dsizeOH [2]; 
    wire[3:0] fragmenter_1__GEN =~ fragmenter_1_dFragnum ; 
    wire[2:0] fragmenter_1_dFirst_size_hi = fragmenter_1_dFragnum [3:1]&{1'h1, fragmenter_1__GEN [3:2]}; 
    wire[3:0] fragmenter_1_dFirst_size_lo ={ fragmenter_1_dFragnum [0], fragmenter_1_dsizeOH1 ,1'h1}&{ fragmenter_1__GEN [1:0],~ fragmenter_1_dsizeOH1 }; 
    wire[3:0] fragmenter_1__dFirst_size_T_8 ={1'h0, fragmenter_1_dFirst_size_hi }| fragmenter_1_dFirst_size_lo ; 
    wire[1:0] fragmenter_1_dFirst_size_hi_1 = fragmenter_1__dFirst_size_T_8 [3:2]; 
    wire[1:0] fragmenter_1_dFirst_size_lo_1 = fragmenter_1__dFirst_size_T_8 [1:0]; 
    wire[2:0] fragmenter_1_dFirst_size ={| fragmenter_1_dFirst_size_hi ,| fragmenter_1_dFirst_size_hi_1 , fragmenter_1_dFirst_size_hi_1 [1]| fragmenter_1_dFirst_size_lo_1 [1]}; 
    wire fragmenter_1_doEarlyAck = fragmenter_1_nodeOut_d_bits_source [5]; 
    wire fragmenter_1_drop =~ fragmenter_1_dHasData &~( fragmenter_1_doEarlyAck  ?  fragmenter_1_dFirst : fragmenter_1_dLast ); 
    wire fragmenter_1_nodeOut_d_ready = fragmenter_1_nodeIn_d_ready | fragmenter_1_drop ; 
    wire fragmenter_1_nodeIn_d_valid = fragmenter_1_nodeOut_d_valid &~ fragmenter_1_drop ; 
    wire[4:0] fragmenter_1_nodeIn_d_bits_source = fragmenter_1_nodeOut_d_bits_source [10:6]; 
    wire[2:0] fragmenter_1_nodeIn_d_bits_size = fragmenter_1_dFirst  ?  fragmenter_1_dFirst_size : fragmenter_1_dOrig ; 
    wire[2:0] fragmenter_1_aFrag = fragmenter_1__repeater_io_deq_bits_size >3'h2 ? 3'h2: fragmenter_1__repeater_io_deq_bits_size ; 
    wire[12:0] fragmenter_1__aOrigOH1_T_1 =13'h3F<< fragmenter_1__repeater_io_deq_bits_size ; 
    wire[5:0] fragmenter_1_aOrigOH1 =~( fragmenter_1__aOrigOH1_T_1 [5:0]); 
    wire[8:0] fragmenter_1__aFragOH1_T_1 =9'h3<< fragmenter_1_aFrag ; 
    wire[1:0] fragmenter_1_aFragOH1 =~( fragmenter_1__aFragOH1_T_1 [1:0]); 
    wire fragmenter_1_aHasData =~( fragmenter_1__repeater_io_deq_bits_opcode [2]); 
    wire[1:0] fragmenter_1_aMask = fragmenter_1_aHasData  ? 2'h0: fragmenter_1_aFragOH1 ; reg[3:0] fragmenter_1_gennum ; 
    wire fragmenter_1_aFirst = fragmenter_1_gennum ==4'h0; 
    wire[3:0] fragmenter_1_old_gennum1 = fragmenter_1_aFirst  ?  fragmenter_1_aOrigOH1 [5:2]: fragmenter_1_gennum -4'h1; 
    wire[3:0] fragmenter_1_new_gennum = fragmenter_1_old_gennum1 ; 
    wire[3:0] fragmenter_1_aFragnum = fragmenter_1_old_gennum1 ; 
    wire fragmenter_1_aLast = fragmenter_1_aFragnum ==4'h0; 
    reg fragmenter_1_aToggle_r ; 
    wire fragmenter_1_aToggle =~( fragmenter_1_aFirst  ?  fragmenter_1_dToggle : fragmenter_1_aToggle_r ); 
    wire fragmenter_1_aFull = fragmenter_1__repeater_io_deq_bits_opcode ==3'h0; 
    wire[31:0] fragmenter_1_nodeOut_a_bits_address ={ fragmenter_1__repeater_io_deq_bits_address [31:6], fragmenter_1__repeater_io_deq_bits_address [5:0]|{~( fragmenter_1_old_gennum1 |~( fragmenter_1_aOrigOH1 [5:2])),2'h0}}; 
    wire[4:0] fragmenter_1_nodeOut_a_bits_source_lo ={ fragmenter_1_aToggle , fragmenter_1_aFragnum }; 
    wire[5:0] fragmenter_1_nodeOut_a_bits_source_hi ={ fragmenter_1__repeater_io_deq_bits_source , fragmenter_1_aFull }; 
    wire[10:0] fragmenter_1_nodeOut_a_bits_source ={ fragmenter_1_nodeOut_a_bits_source_hi , fragmenter_1_nodeOut_a_bits_source_lo }; 
    wire[1:0] fragmenter_1_nodeOut_a_bits_size = fragmenter_1_aFrag [1:0]; 
  always @( posedge  fragmenter_1_clock )
         begin 
             if (~ fragmenter_1_reset &~(~ fragmenter_1__repeater_io_full |~ fragmenter_1_aHasData ))
                 begin 
                     if (1)$error("Assertion failed\n    at Fragmenter.scala:311 assert (!repeater.io.full || !aHasData)\n");
                     if (1)$fatal;
                 end 
             if (~ fragmenter_1_reset &~(~ fragmenter_1__repeater_io_full |(& fragmenter_1__repeater_io_deq_bits_mask )))
                 begin 
                     if (1)$error("Assertion failed\n    at Fragmenter.scala:314 assert (!repeater.io.full || in_a.bits.mask === fullMask)\n");
                     if (1)$fatal;
                 end 
         end
    wire[3:0] fragmenter_1_nodeOut_a_bits_mask = fragmenter_1__repeater_io_full  ? 4'hF: fragmenter_1_nodeIn_a_bits_mask ; 
    wire fragmenter_1_nodeOut_a_valid ; 
    wire fragmenter_1__GEN_0 = fragmenter_1_nodeOut_d_ready & fragmenter_1_nodeOut_d_valid ; 
    wire fragmenter_1__GEN_1 = fragmenter_1__GEN_0 & fragmenter_1_dFirst ; 
  always @( posedge  fragmenter_1_clock )
         begin 
             if ( fragmenter_1_reset )
                 begin  
                     fragmenter_1_acknum  <=4'h0; 
                     fragmenter_1_dToggle  <=1'h0; 
                     fragmenter_1_gennum  <=4'h0;
                 end 
              else 
                 begin 
                     if ( fragmenter_1__GEN_0 )
                         begin 
                             if ( fragmenter_1_dFirst ) 
                                 fragmenter_1_acknum  <= fragmenter_1_dFirst_acknum ;
                              else  
                                 fragmenter_1_acknum  <= fragmenter_1_acknum -{3'h0, fragmenter_1_ack_decrement };
                         end 
                     if ( fragmenter_1__GEN_1 ) 
                         fragmenter_1_dToggle  <= fragmenter_1_nodeOut_d_bits_source [4];
                     if ( fragmenter_1_nodeOut_a_ready & fragmenter_1_nodeOut_a_valid ) 
                         fragmenter_1_gennum  <= fragmenter_1_new_gennum ;
                 end 
             if ( fragmenter_1__GEN_1 ) 
                 fragmenter_1_dOrig  <= fragmenter_1_dFirst_size ;
             if ( fragmenter_1_aFirst ) 
                 fragmenter_1_aToggle_r  <= fragmenter_1_dToggle ;
         end
    wire fragmenter_1_repeater_clock;
    wire fragmenter_1_repeater_reset;
    wire fragmenter_1_repeater_io_repeat;
    wire fragmenter_1_repeater_io_full;
    wire fragmenter_1_repeater_io_enq_ready;
    wire fragmenter_1_repeater_io_enq_valid;
    wire[2:0] fragmenter_1_repeater_io_enq_bits_opcode;
    wire[2:0] fragmenter_1_repeater_io_enq_bits_param;
    wire[2:0] fragmenter_1_repeater_io_enq_bits_size;
    wire[4:0] fragmenter_1_repeater_io_enq_bits_source;
    wire[31:0] fragmenter_1_repeater_io_enq_bits_address;
    wire[3:0] fragmenter_1_repeater_io_enq_bits_mask;
    wire[31:0] fragmenter_1_repeater_io_enq_bits_data;
    wire fragmenter_1_repeater_io_enq_bits_corrupt;
    wire fragmenter_1_repeater_io_deq_ready;
    wire fragmenter_1_repeater_io_deq_valid;
    wire[2:0] fragmenter_1_repeater_io_deq_bits_opcode;
    wire[2:0] fragmenter_1_repeater_io_deq_bits_param;
    wire[2:0] fragmenter_1_repeater_io_deq_bits_size;
    wire[4:0] fragmenter_1_repeater_io_deq_bits_source;
    wire[31:0] fragmenter_1_repeater_io_deq_bits_address;
    wire[3:0] fragmenter_1_repeater_io_deq_bits_mask;
    wire fragmenter_1_repeater_io_deq_bits_corrupt;

    reg fragmenter_1_repeater_full ; reg[2:0] fragmenter_1_repeater_saved_opcode ; reg[2:0] fragmenter_1_repeater_saved_param ; reg[2:0] fragmenter_1_repeater_saved_size ; reg[4:0] fragmenter_1_repeater_saved_source ; reg[31:0] fragmenter_1_repeater_saved_address ; reg[3:0] fragmenter_1_repeater_saved_mask ; reg[31:0] fragmenter_1_repeater_saved_data ; 
    reg fragmenter_1_repeater_saved_corrupt ; 
    wire fragmenter_1_repeater__io_deq_valid_output = fragmenter_1_repeater_io_enq_valid | fragmenter_1_repeater_full ; 
    wire fragmenter_1_repeater__io_enq_ready_output = fragmenter_1_repeater_io_deq_ready &~ fragmenter_1_repeater_full ; 
    wire fragmenter_1_repeater__GEN = fragmenter_1_repeater__io_enq_ready_output & fragmenter_1_repeater_io_enq_valid & fragmenter_1_repeater_io_repeat ; 
  always @( posedge  fragmenter_1_repeater_clock )
         begin 
             if ( fragmenter_1_repeater_reset ) 
                 fragmenter_1_repeater_full  <=1'h0;
              else  
                 fragmenter_1_repeater_full  <=~( fragmenter_1_repeater_io_deq_ready & fragmenter_1_repeater__io_deq_valid_output &~ fragmenter_1_repeater_io_repeat )&( fragmenter_1_repeater__GEN | fragmenter_1_repeater_full );
             if ( fragmenter_1_repeater__GEN )
                 begin  
                     fragmenter_1_repeater_saved_opcode  <= fragmenter_1_repeater_io_enq_bits_opcode ; 
                     fragmenter_1_repeater_saved_param  <= fragmenter_1_repeater_io_enq_bits_param ; 
                     fragmenter_1_repeater_saved_size  <= fragmenter_1_repeater_io_enq_bits_size ; 
                     fragmenter_1_repeater_saved_source  <= fragmenter_1_repeater_io_enq_bits_source ; 
                     fragmenter_1_repeater_saved_address  <= fragmenter_1_repeater_io_enq_bits_address ; 
                     fragmenter_1_repeater_saved_mask  <= fragmenter_1_repeater_io_enq_bits_mask ; 
                     fragmenter_1_repeater_saved_data  <= fragmenter_1_repeater_io_enq_bits_data ; 
                     fragmenter_1_repeater_saved_corrupt  <= fragmenter_1_repeater_io_enq_bits_corrupt ;
                 end 
         end
  assign  fragmenter_1_repeater_io_full = fragmenter_1_repeater_full ; 
  assign  fragmenter_1_repeater_io_enq_ready = fragmenter_1_repeater__io_enq_ready_output ; 
  assign  fragmenter_1_repeater_io_deq_valid = fragmenter_1_repeater__io_deq_valid_output ; 
  assign  fragmenter_1_repeater_io_deq_bits_opcode = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_opcode : fragmenter_1_repeater_io_enq_bits_opcode ; 
  assign  fragmenter_1_repeater_io_deq_bits_param = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_param : fragmenter_1_repeater_io_enq_bits_param ; 
  assign  fragmenter_1_repeater_io_deq_bits_size = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_size : fragmenter_1_repeater_io_enq_bits_size ; 
  assign  fragmenter_1_repeater_io_deq_bits_source = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_source : fragmenter_1_repeater_io_enq_bits_source ; 
  assign  fragmenter_1_repeater_io_deq_bits_address = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_address : fragmenter_1_repeater_io_enq_bits_address ; 
  assign  fragmenter_1_repeater_io_deq_bits_mask = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_mask : fragmenter_1_repeater_io_enq_bits_mask ; 
  assign  fragmenter_1_repeater_io_deq_bits_corrupt = fragmenter_1_repeater_full  ?  fragmenter_1_repeater_saved_corrupt : fragmenter_1_repeater_io_enq_bits_corrupt ;
    assign fragmenter_1_repeater_clock = fragmenter_1_clock;
    assign fragmenter_1_repeater_reset = fragmenter_1_reset;
    assign fragmenter_1_repeater_io_repeat = ~fragmenter_1_aHasData&(|fragmenter_1_aFragnum);
    assign fragmenter_1__repeater_io_full = fragmenter_1_repeater_io_full;
    assign fragmenter_1_nodeIn_a_ready = fragmenter_1_repeater_io_enq_ready;
    assign fragmenter_1_repeater_io_enq_valid = fragmenter_1_nodeIn_a_valid;
    assign fragmenter_1_repeater_io_enq_bits_opcode = fragmenter_1_nodeIn_a_bits_opcode;
    assign fragmenter_1_repeater_io_enq_bits_param = fragmenter_1_nodeIn_a_bits_param;
    assign fragmenter_1_repeater_io_enq_bits_size = fragmenter_1_nodeIn_a_bits_size;
    assign fragmenter_1_repeater_io_enq_bits_source = fragmenter_1_nodeIn_a_bits_source;
    assign fragmenter_1_repeater_io_enq_bits_address = fragmenter_1_nodeIn_a_bits_address;
    assign fragmenter_1_repeater_io_enq_bits_mask = fragmenter_1_nodeIn_a_bits_mask;
    assign fragmenter_1_repeater_io_enq_bits_data = fragmenter_1_nodeIn_a_bits_data;
    assign fragmenter_1_repeater_io_enq_bits_corrupt = fragmenter_1_nodeIn_a_bits_corrupt;
    assign fragmenter_1_repeater_io_deq_ready = fragmenter_1_nodeOut_a_ready;
    assign fragmenter_1_nodeOut_a_valid = fragmenter_1_repeater_io_deq_valid;
    assign fragmenter_1__repeater_io_deq_bits_opcode = fragmenter_1_repeater_io_deq_bits_opcode;
    assign fragmenter_1_nodeOut_a_bits_param = fragmenter_1_repeater_io_deq_bits_param;
    assign fragmenter_1__repeater_io_deq_bits_size = fragmenter_1_repeater_io_deq_bits_size;
    assign fragmenter_1__repeater_io_deq_bits_source = fragmenter_1_repeater_io_deq_bits_source;
    assign fragmenter_1__repeater_io_deq_bits_address = fragmenter_1_repeater_io_deq_bits_address;
    assign fragmenter_1__repeater_io_deq_bits_mask = fragmenter_1_repeater_io_deq_bits_mask;
    assign fragmenter_1_nodeOut_a_bits_corrupt = fragmenter_1_repeater_io_deq_bits_corrupt;
     
    wire[2:0] fragmenter_1_nodeOut_a_bits_opcode ; 
  assign  fragmenter_1_nodeOut_a_bits_opcode = fragmenter_1__repeater_io_deq_bits_opcode ; 
  assign  fragmenter_1_auto_in_a_ready = fragmenter_1_nodeIn_a_ready ; 
  assign  fragmenter_1_auto_in_d_valid = fragmenter_1_nodeIn_d_valid ; 
  assign  fragmenter_1_auto_in_d_bits_opcode = fragmenter_1_nodeIn_d_bits_opcode ; 
  assign  fragmenter_1_auto_in_d_bits_size = fragmenter_1_nodeIn_d_bits_size ; 
  assign  fragmenter_1_auto_in_d_bits_source = fragmenter_1_nodeIn_d_bits_source ; 
  assign  fragmenter_1_auto_in_d_bits_data = fragmenter_1_nodeIn_d_bits_data ; 
  assign  fragmenter_1_auto_out_a_valid = fragmenter_1_nodeOut_a_valid ; 
  assign  fragmenter_1_auto_out_a_bits_opcode = fragmenter_1_nodeOut_a_bits_opcode ; 
  assign  fragmenter_1_auto_out_a_bits_param = fragmenter_1_nodeOut_a_bits_param ; 
  assign  fragmenter_1_auto_out_a_bits_size = fragmenter_1_nodeOut_a_bits_size ; 
  assign  fragmenter_1_auto_out_a_bits_source = fragmenter_1_nodeOut_a_bits_source ; 
  assign  fragmenter_1_auto_out_a_bits_address = fragmenter_1_nodeOut_a_bits_address ; 
  assign  fragmenter_1_auto_out_a_bits_mask = fragmenter_1_nodeOut_a_bits_mask ; 
  assign  fragmenter_1_auto_out_a_bits_data = fragmenter_1_nodeOut_a_bits_data ; 
  assign  fragmenter_1_auto_out_a_bits_corrupt = fragmenter_1_nodeOut_a_bits_corrupt ; 
  assign  fragmenter_1_auto_out_d_ready = fragmenter_1_nodeOut_d_ready ;
    assign fragmenter_1_clock = clock;
    assign fragmenter_1_reset = reset;
    assign tlSlaveXbar_nodeOut_a_ready = fragmenter_1_auto_in_a_ready;
    assign fragmenter_1_auto_in_a_valid = tlSlaveXbar_nodeOut_a_valid;
    assign fragmenter_1_auto_in_a_bits_opcode = tlSlaveXbar_nodeOut_a_bits_opcode;
    assign fragmenter_1_auto_in_a_bits_param = tlSlaveXbar_nodeOut_a_bits_param;
    assign fragmenter_1_auto_in_a_bits_size = tlSlaveXbar_nodeOut_a_bits_size;
    assign fragmenter_1_auto_in_a_bits_source = tlSlaveXbar_nodeOut_a_bits_source;
    assign fragmenter_1_auto_in_a_bits_address = tlSlaveXbar_nodeOut_a_bits_address;
    assign fragmenter_1_auto_in_a_bits_mask = tlSlaveXbar_nodeOut_a_bits_mask;
    assign fragmenter_1_auto_in_a_bits_data = tlSlaveXbar_nodeOut_a_bits_data;
    assign fragmenter_1_auto_in_a_bits_corrupt = tlSlaveXbar_nodeOut_a_bits_corrupt;
    assign fragmenter_1_auto_in_d_ready = tlSlaveXbar_nodeOut_d_ready;
    assign tlSlaveXbar_nodeOut_d_valid = fragmenter_1_auto_in_d_valid;
    assign tlSlaveXbar_nodeOut_d_bits_opcode = fragmenter_1_auto_in_d_bits_opcode;
    assign tlSlaveXbar_nodeOut_d_bits_size = fragmenter_1_auto_in_d_bits_size;
    assign tlSlaveXbar_nodeOut_d_bits_source = fragmenter_1_auto_in_d_bits_source;
    assign tlSlaveXbar_nodeOut_d_bits_data = fragmenter_1_auto_in_d_bits_data;
    assign fragmenter_1_auto_out_a_ready = _dtim_adapter_auto_in_a_ready;
    assign _fragmenter_1_auto_out_a_valid = fragmenter_1_auto_out_a_valid;
    assign _fragmenter_1_auto_out_a_bits_opcode = fragmenter_1_auto_out_a_bits_opcode;
    assign _fragmenter_1_auto_out_a_bits_param = fragmenter_1_auto_out_a_bits_param;
    assign _fragmenter_1_auto_out_a_bits_size = fragmenter_1_auto_out_a_bits_size;
    assign _fragmenter_1_auto_out_a_bits_source = fragmenter_1_auto_out_a_bits_source;
    assign _fragmenter_1_auto_out_a_bits_address = fragmenter_1_auto_out_a_bits_address;
    assign _fragmenter_1_auto_out_a_bits_mask = fragmenter_1_auto_out_a_bits_mask;
    assign _fragmenter_1_auto_out_a_bits_data = fragmenter_1_auto_out_a_bits_data;
    assign _fragmenter_1_auto_out_a_bits_corrupt = fragmenter_1_auto_out_a_bits_corrupt;
    assign _fragmenter_1_auto_out_d_ready = fragmenter_1_auto_out_d_ready;
    assign fragmenter_1_auto_out_d_valid = _dtim_adapter_auto_in_d_valid;
    assign fragmenter_1_auto_out_d_bits_opcode = _dtim_adapter_auto_in_d_bits_opcode;
    assign fragmenter_1_auto_out_d_bits_size = _dtim_adapter_auto_in_d_bits_size;
    assign fragmenter_1_auto_out_d_bits_source = _dtim_adapter_auto_in_d_bits_source;
    assign fragmenter_1_auto_out_d_bits_data = _dtim_adapter_auto_in_d_bits_data;
    
  wire dcacheArb_clock;
    wire dcacheArb_io_requestor_0_req_ready;
    wire dcacheArb_io_requestor_0_req_valid;
    wire[31:0] dcacheArb_io_requestor_0_req_bits_addr;
    wire[6:0] dcacheArb_io_requestor_0_req_bits_tag;
    wire[4:0] dcacheArb_io_requestor_0_req_bits_cmd;
    wire[1:0] dcacheArb_io_requestor_0_req_bits_size;
    wire dcacheArb_io_requestor_0_req_bits_signed;
    wire dcacheArb_io_requestor_0_req_bits_dv;
    wire dcacheArb_io_requestor_0_s1_kill;
    wire[31:0] dcacheArb_io_requestor_0_s1_data_data;
    wire dcacheArb_io_requestor_0_s2_nack;
    wire dcacheArb_io_requestor_0_resp_valid;
    wire[6:0] dcacheArb_io_requestor_0_resp_bits_tag;
    wire[31:0] dcacheArb_io_requestor_0_resp_bits_data;
    wire dcacheArb_io_requestor_0_resp_bits_replay;
    wire dcacheArb_io_requestor_0_resp_bits_has_data;
    wire[31:0] dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
    wire dcacheArb_io_requestor_0_replay_next;
    wire dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_ma_st;
    wire dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_pf_st;
    wire dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_ae_st;
    wire dcacheArb_io_requestor_0_ordered;
    wire dcacheArb_io_requestor_0_perf_grant;
    wire dcacheArb_io_requestor_1_req_ready;
    wire dcacheArb_io_requestor_1_req_valid;
    wire[31:0] dcacheArb_io_requestor_1_req_bits_addr;
    wire[4:0] dcacheArb_io_requestor_1_req_bits_cmd;
    wire[1:0] dcacheArb_io_requestor_1_req_bits_size;
    wire dcacheArb_io_requestor_1_s1_kill;
    wire[31:0] dcacheArb_io_requestor_1_s1_data_data;
    wire[3:0] dcacheArb_io_requestor_1_s1_data_mask;
    wire dcacheArb_io_requestor_1_s2_nack;
    wire dcacheArb_io_requestor_1_resp_valid;
    wire[31:0] dcacheArb_io_requestor_1_resp_bits_data_raw;
    wire dcacheArb_io_mem_req_ready;
    wire dcacheArb_io_mem_req_valid;
    wire[31:0] dcacheArb_io_mem_req_bits_addr;
    wire[6:0] dcacheArb_io_mem_req_bits_tag;
    wire[4:0] dcacheArb_io_mem_req_bits_cmd;
    wire[1:0] dcacheArb_io_mem_req_bits_size;
    wire dcacheArb_io_mem_req_bits_signed;
    wire[1:0] dcacheArb_io_mem_req_bits_dprv;
    wire dcacheArb_io_mem_req_bits_dv;
    wire dcacheArb_io_mem_req_bits_phys;
    wire dcacheArb_io_mem_req_bits_no_xcpt;
    wire dcacheArb_io_mem_s1_kill;
    wire[31:0] dcacheArb_io_mem_s1_data_data;
    wire[3:0] dcacheArb_io_mem_s1_data_mask;
    wire dcacheArb_io_mem_s2_nack;
    wire dcacheArb_io_mem_resp_valid;
    wire[6:0] dcacheArb_io_mem_resp_bits_tag;
    wire[31:0] dcacheArb_io_mem_resp_bits_data;
    wire dcacheArb_io_mem_resp_bits_replay;
    wire dcacheArb_io_mem_resp_bits_has_data;
    wire[31:0] dcacheArb_io_mem_resp_bits_data_word_bypass;
    wire[31:0] dcacheArb_io_mem_resp_bits_data_raw;
    wire dcacheArb_io_mem_replay_next;
    wire dcacheArb_io_mem_s2_xcpt_ma_ld;
    wire dcacheArb_io_mem_s2_xcpt_ma_st;
    wire dcacheArb_io_mem_s2_xcpt_pf_ld;
    wire dcacheArb_io_mem_s2_xcpt_pf_st;
    wire dcacheArb_io_mem_s2_xcpt_ae_ld;
    wire dcacheArb_io_mem_s2_xcpt_ae_st;
    wire dcacheArb_io_mem_ordered;
    wire dcacheArb_io_mem_perf_grant;

    reg dcacheArb_s1_id ; 
    reg dcacheArb_s2_id ; 
    wire dcacheArb_tag_hit_1 = dcacheArb_io_mem_resp_bits_tag [0]; 
    wire dcacheArb_tag_hit =~ dcacheArb_tag_hit_1 ; 
  always @( posedge  dcacheArb_clock )
         begin  
             dcacheArb_s1_id  <=~ dcacheArb_io_requestor_0_req_valid ; 
             dcacheArb_s2_id  <= dcacheArb_s1_id ;
         end
  assign  dcacheArb_io_requestor_0_req_ready = dcacheArb_io_mem_req_ready ; 
  assign  dcacheArb_io_requestor_0_s2_nack = dcacheArb_io_mem_s2_nack &~ dcacheArb_s2_id ; 
  assign  dcacheArb_io_requestor_0_resp_valid = dcacheArb_io_mem_resp_valid & dcacheArb_tag_hit ; 
  assign  dcacheArb_io_requestor_0_resp_bits_tag ={1'h0, dcacheArb_io_mem_resp_bits_tag [6:1]}; 
  assign  dcacheArb_io_requestor_0_resp_bits_data = dcacheArb_io_mem_resp_bits_data ; 
  assign  dcacheArb_io_requestor_0_resp_bits_replay = dcacheArb_io_mem_resp_bits_replay ; 
  assign  dcacheArb_io_requestor_0_resp_bits_has_data = dcacheArb_io_mem_resp_bits_has_data ; 
  assign  dcacheArb_io_requestor_0_resp_bits_data_word_bypass = dcacheArb_io_mem_resp_bits_data_word_bypass ; 
  assign  dcacheArb_io_requestor_0_replay_next = dcacheArb_io_mem_replay_next ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ma_ld = dcacheArb_io_mem_s2_xcpt_ma_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ma_st = dcacheArb_io_mem_s2_xcpt_ma_st ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_pf_ld = dcacheArb_io_mem_s2_xcpt_pf_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_pf_st = dcacheArb_io_mem_s2_xcpt_pf_st ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ae_ld = dcacheArb_io_mem_s2_xcpt_ae_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ae_st = dcacheArb_io_mem_s2_xcpt_ae_st ; 
  assign  dcacheArb_io_requestor_0_ordered = dcacheArb_io_mem_ordered ; 
  assign  dcacheArb_io_requestor_0_perf_grant = dcacheArb_io_mem_perf_grant ; 
  assign  dcacheArb_io_requestor_1_req_ready = dcacheArb_io_mem_req_ready &~ dcacheArb_io_requestor_0_req_valid ; 
  assign  dcacheArb_io_requestor_1_s2_nack = dcacheArb_io_mem_s2_nack & dcacheArb_s2_id ; 
  assign  dcacheArb_io_requestor_1_resp_valid = dcacheArb_io_mem_resp_valid & dcacheArb_tag_hit_1 ; 
  assign  dcacheArb_io_requestor_1_resp_bits_data_raw = dcacheArb_io_mem_resp_bits_data_raw ; 
  assign  dcacheArb_io_mem_req_valid = dcacheArb_io_requestor_0_req_valid | dcacheArb_io_requestor_1_req_valid ; 
  assign  dcacheArb_io_mem_req_bits_addr = dcacheArb_io_requestor_0_req_valid  ?  dcacheArb_io_requestor_0_req_bits_addr : dcacheArb_io_requestor_1_req_bits_addr ; 
  assign  dcacheArb_io_mem_req_bits_tag = dcacheArb_io_requestor_0_req_valid  ? { dcacheArb_io_requestor_0_req_bits_tag [5:0],1'h0}:7'h1; 
  assign  dcacheArb_io_mem_req_bits_cmd = dcacheArb_io_requestor_0_req_valid  ?  dcacheArb_io_requestor_0_req_bits_cmd : dcacheArb_io_requestor_1_req_bits_cmd ; 
  assign  dcacheArb_io_mem_req_bits_size = dcacheArb_io_requestor_0_req_valid  ?  dcacheArb_io_requestor_0_req_bits_size : dcacheArb_io_requestor_1_req_bits_size ; 
  assign  dcacheArb_io_mem_req_bits_signed = dcacheArb_io_requestor_0_req_valid & dcacheArb_io_requestor_0_req_bits_signed ; 
  assign  dcacheArb_io_mem_req_bits_dprv ={2{ dcacheArb_io_requestor_0_req_valid }}; 
  assign  dcacheArb_io_mem_req_bits_dv = dcacheArb_io_requestor_0_req_valid & dcacheArb_io_requestor_0_req_bits_dv ; 
  assign  dcacheArb_io_mem_req_bits_phys =~ dcacheArb_io_requestor_0_req_valid ; 
  assign  dcacheArb_io_mem_req_bits_no_xcpt =~ dcacheArb_io_requestor_0_req_valid ; 
  assign  dcacheArb_io_mem_s1_kill = dcacheArb_s1_id  ?  dcacheArb_io_requestor_1_s1_kill : dcacheArb_io_requestor_0_s1_kill ; 
  assign  dcacheArb_io_mem_s1_data_data = dcacheArb_s1_id  ?  dcacheArb_io_requestor_1_s1_data_data : dcacheArb_io_requestor_0_s1_data_data ; 
  assign  dcacheArb_io_mem_s1_data_mask = dcacheArb_s1_id  ?  dcacheArb_io_requestor_1_s1_data_mask :4'h0;
    assign dcacheArb_clock = clock;
    assign _dcacheArb_io_requestor_0_req_ready = dcacheArb_io_requestor_0_req_ready;
    assign dcacheArb_io_requestor_0_req_valid = _core_io_dmem_req_valid;
    assign dcacheArb_io_requestor_0_req_bits_addr = _core_io_dmem_req_bits_addr;
    assign dcacheArb_io_requestor_0_req_bits_tag = _core_io_dmem_req_bits_tag;
    assign dcacheArb_io_requestor_0_req_bits_cmd = _core_io_dmem_req_bits_cmd;
    assign dcacheArb_io_requestor_0_req_bits_size = _core_io_dmem_req_bits_size;
    assign dcacheArb_io_requestor_0_req_bits_signed = _core_io_dmem_req_bits_signed;
    assign dcacheArb_io_requestor_0_req_bits_dv = _core_io_dmem_req_bits_dv;
    assign dcacheArb_io_requestor_0_s1_kill = _core_io_dmem_s1_kill;
    assign dcacheArb_io_requestor_0_s1_data_data = _core_io_dmem_s1_data_data;
    assign _dcacheArb_io_requestor_0_s2_nack = dcacheArb_io_requestor_0_s2_nack;
    assign _dcacheArb_io_requestor_0_resp_valid = dcacheArb_io_requestor_0_resp_valid;
    assign _dcacheArb_io_requestor_0_resp_bits_tag = dcacheArb_io_requestor_0_resp_bits_tag;
    assign _dcacheArb_io_requestor_0_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data;
    assign _dcacheArb_io_requestor_0_resp_bits_replay = dcacheArb_io_requestor_0_resp_bits_replay;
    assign _dcacheArb_io_requestor_0_resp_bits_has_data = dcacheArb_io_requestor_0_resp_bits_has_data;
    assign _dcacheArb_io_requestor_0_resp_bits_data_word_bypass = dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
    assign _dcacheArb_io_requestor_0_replay_next = dcacheArb_io_requestor_0_replay_next;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ma_ld = dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ma_st = dcacheArb_io_requestor_0_s2_xcpt_ma_st;
    assign _dcacheArb_io_requestor_0_s2_xcpt_pf_ld = dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_pf_st = dcacheArb_io_requestor_0_s2_xcpt_pf_st;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ae_st = dcacheArb_io_requestor_0_s2_xcpt_ae_st;
    assign _dcacheArb_io_requestor_0_ordered = dcacheArb_io_requestor_0_ordered;
    assign _dcacheArb_io_requestor_0_perf_grant = dcacheArb_io_requestor_0_perf_grant;
    assign _dcacheArb_io_requestor_1_req_ready = dcacheArb_io_requestor_1_req_ready;
    assign dcacheArb_io_requestor_1_req_valid = _dtim_adapter_io_dmem_req_valid;
    assign dcacheArb_io_requestor_1_req_bits_addr = _dtim_adapter_io_dmem_req_bits_addr;
    assign dcacheArb_io_requestor_1_req_bits_cmd = _dtim_adapter_io_dmem_req_bits_cmd;
    assign dcacheArb_io_requestor_1_req_bits_size = _dtim_adapter_io_dmem_req_bits_size;
    assign dcacheArb_io_requestor_1_s1_kill = _dtim_adapter_io_dmem_s1_kill;
    assign dcacheArb_io_requestor_1_s1_data_data = _dtim_adapter_io_dmem_s1_data_data;
    assign dcacheArb_io_requestor_1_s1_data_mask = _dtim_adapter_io_dmem_s1_data_mask;
    assign _dcacheArb_io_requestor_1_s2_nack = dcacheArb_io_requestor_1_s2_nack;
    assign _dcacheArb_io_requestor_1_resp_valid = dcacheArb_io_requestor_1_resp_valid;
    assign _dcacheArb_io_requestor_1_resp_bits_data_raw = dcacheArb_io_requestor_1_resp_bits_data_raw;
    assign dcacheArb_io_mem_req_ready = _dcache_io_cpu_req_ready;
    assign _dcacheArb_io_mem_req_valid = dcacheArb_io_mem_req_valid;
    assign _dcacheArb_io_mem_req_bits_addr = dcacheArb_io_mem_req_bits_addr;
    assign _dcacheArb_io_mem_req_bits_tag = dcacheArb_io_mem_req_bits_tag;
    assign _dcacheArb_io_mem_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd;
    assign _dcacheArb_io_mem_req_bits_size = dcacheArb_io_mem_req_bits_size;
    assign _dcacheArb_io_mem_req_bits_signed = dcacheArb_io_mem_req_bits_signed;
    assign _dcacheArb_io_mem_req_bits_dprv = dcacheArb_io_mem_req_bits_dprv;
    assign _dcacheArb_io_mem_req_bits_dv = dcacheArb_io_mem_req_bits_dv;
    assign _dcacheArb_io_mem_req_bits_phys = dcacheArb_io_mem_req_bits_phys;
    assign _dcacheArb_io_mem_req_bits_no_xcpt = dcacheArb_io_mem_req_bits_no_xcpt;
    assign _dcacheArb_io_mem_s1_kill = dcacheArb_io_mem_s1_kill;
    assign _dcacheArb_io_mem_s1_data_data = dcacheArb_io_mem_s1_data_data;
    assign _dcacheArb_io_mem_s1_data_mask = dcacheArb_io_mem_s1_data_mask;
    assign dcacheArb_io_mem_s2_nack = _dcache_io_cpu_s2_nack;
    assign dcacheArb_io_mem_resp_valid = _dcache_io_cpu_resp_valid;
    assign dcacheArb_io_mem_resp_bits_tag = _dcache_io_cpu_resp_bits_tag;
    assign dcacheArb_io_mem_resp_bits_data = _dcache_io_cpu_resp_bits_data;
    assign dcacheArb_io_mem_resp_bits_replay = _dcache_io_cpu_resp_bits_replay;
    assign dcacheArb_io_mem_resp_bits_has_data = _dcache_io_cpu_resp_bits_has_data;
    assign dcacheArb_io_mem_resp_bits_data_word_bypass = _dcache_io_cpu_resp_bits_data_word_bypass;
    assign dcacheArb_io_mem_resp_bits_data_raw = _dcache_io_cpu_resp_bits_data_raw;
    assign dcacheArb_io_mem_replay_next = _dcache_io_cpu_replay_next;
    assign dcacheArb_io_mem_s2_xcpt_ma_ld = _dcache_io_cpu_s2_xcpt_ma_ld;
    assign dcacheArb_io_mem_s2_xcpt_ma_st = _dcache_io_cpu_s2_xcpt_ma_st;
    assign dcacheArb_io_mem_s2_xcpt_pf_ld = _dcache_io_cpu_s2_xcpt_pf_ld;
    assign dcacheArb_io_mem_s2_xcpt_pf_st = _dcache_io_cpu_s2_xcpt_pf_st;
    assign dcacheArb_io_mem_s2_xcpt_ae_ld = _dcache_io_cpu_s2_xcpt_ae_ld;
    assign dcacheArb_io_mem_s2_xcpt_ae_st = _dcache_io_cpu_s2_xcpt_ae_st;
    assign dcacheArb_io_mem_ordered = _dcache_io_cpu_ordered;
    assign dcacheArb_io_mem_perf_grant = _dcache_io_cpu_perf_grant;
    
  wire ptw_clock;
    wire ptw_reset;
    wire[19:0] ptw_io_requestor_0_req_bits_bits_addr;
    wire ptw_io_requestor_0_req_bits_bits_need_gpa;
    wire ptw_io_requestor_0_req_bits_bits_vstage1;
    wire ptw_io_requestor_0_req_bits_bits_stage2;
    wire ptw_io_requestor_0_resp_bits_ae_ptw;
    wire ptw_io_requestor_0_resp_bits_ae_final;
    wire ptw_io_requestor_0_resp_bits_pf;
    wire ptw_io_requestor_0_resp_bits_gf;
    wire ptw_io_requestor_0_resp_bits_hr;
    wire ptw_io_requestor_0_resp_bits_hw;
    wire ptw_io_requestor_0_resp_bits_hx;
    wire[43:0] ptw_io_requestor_0_resp_bits_pte_ppn;
    wire ptw_io_requestor_0_resp_bits_pte_d;
    wire ptw_io_requestor_0_resp_bits_pte_a;
    wire ptw_io_requestor_0_resp_bits_pte_g;
    wire ptw_io_requestor_0_resp_bits_pte_u;
    wire ptw_io_requestor_0_resp_bits_pte_x;
    wire ptw_io_requestor_0_resp_bits_pte_w;
    wire ptw_io_requestor_0_resp_bits_pte_r;
    wire ptw_io_requestor_0_resp_bits_pte_v;
    wire ptw_io_requestor_0_resp_bits_gpa_is_pte;
    wire ptw_io_requestor_0_status_debug;
    wire ptw_io_requestor_0_pmp_0_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_0_cfg_a;
    wire ptw_io_requestor_0_pmp_0_cfg_x;
    wire ptw_io_requestor_0_pmp_0_cfg_w;
    wire ptw_io_requestor_0_pmp_0_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_0_addr;
    wire[31:0] ptw_io_requestor_0_pmp_0_mask;
    wire ptw_io_requestor_0_pmp_1_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_1_cfg_a;
    wire ptw_io_requestor_0_pmp_1_cfg_x;
    wire ptw_io_requestor_0_pmp_1_cfg_w;
    wire ptw_io_requestor_0_pmp_1_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_1_addr;
    wire[31:0] ptw_io_requestor_0_pmp_1_mask;
    wire ptw_io_requestor_0_pmp_2_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_2_cfg_a;
    wire ptw_io_requestor_0_pmp_2_cfg_x;
    wire ptw_io_requestor_0_pmp_2_cfg_w;
    wire ptw_io_requestor_0_pmp_2_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_2_addr;
    wire[31:0] ptw_io_requestor_0_pmp_2_mask;
    wire ptw_io_requestor_0_pmp_3_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_3_cfg_a;
    wire ptw_io_requestor_0_pmp_3_cfg_x;
    wire ptw_io_requestor_0_pmp_3_cfg_w;
    wire ptw_io_requestor_0_pmp_3_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_3_addr;
    wire[31:0] ptw_io_requestor_0_pmp_3_mask;
    wire ptw_io_requestor_0_pmp_4_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_4_cfg_a;
    wire ptw_io_requestor_0_pmp_4_cfg_x;
    wire ptw_io_requestor_0_pmp_4_cfg_w;
    wire ptw_io_requestor_0_pmp_4_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_4_addr;
    wire[31:0] ptw_io_requestor_0_pmp_4_mask;
    wire ptw_io_requestor_0_pmp_5_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_5_cfg_a;
    wire ptw_io_requestor_0_pmp_5_cfg_x;
    wire ptw_io_requestor_0_pmp_5_cfg_w;
    wire ptw_io_requestor_0_pmp_5_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_5_addr;
    wire[31:0] ptw_io_requestor_0_pmp_5_mask;
    wire ptw_io_requestor_0_pmp_6_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_6_cfg_a;
    wire ptw_io_requestor_0_pmp_6_cfg_x;
    wire ptw_io_requestor_0_pmp_6_cfg_w;
    wire ptw_io_requestor_0_pmp_6_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_6_addr;
    wire[31:0] ptw_io_requestor_0_pmp_6_mask;
    wire ptw_io_requestor_0_pmp_7_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_7_cfg_a;
    wire ptw_io_requestor_0_pmp_7_cfg_x;
    wire ptw_io_requestor_0_pmp_7_cfg_w;
    wire ptw_io_requestor_0_pmp_7_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_7_addr;
    wire[31:0] ptw_io_requestor_0_pmp_7_mask;
    wire ptw_io_requestor_1_req_bits_valid;
    wire[19:0] ptw_io_requestor_1_req_bits_bits_addr;
    wire ptw_io_requestor_1_req_bits_bits_need_gpa;
    wire ptw_io_requestor_1_req_bits_bits_vstage1;
    wire ptw_io_requestor_1_req_bits_bits_stage2;
    wire ptw_io_requestor_1_resp_bits_ae_ptw;
    wire ptw_io_requestor_1_resp_bits_ae_final;
    wire ptw_io_requestor_1_resp_bits_pf;
    wire ptw_io_requestor_1_resp_bits_gf;
    wire ptw_io_requestor_1_resp_bits_hr;
    wire ptw_io_requestor_1_resp_bits_hw;
    wire ptw_io_requestor_1_resp_bits_hx;
    wire[43:0] ptw_io_requestor_1_resp_bits_pte_ppn;
    wire ptw_io_requestor_1_resp_bits_pte_d;
    wire ptw_io_requestor_1_resp_bits_pte_a;
    wire ptw_io_requestor_1_resp_bits_pte_g;
    wire ptw_io_requestor_1_resp_bits_pte_u;
    wire ptw_io_requestor_1_resp_bits_pte_x;
    wire ptw_io_requestor_1_resp_bits_pte_w;
    wire ptw_io_requestor_1_resp_bits_pte_r;
    wire ptw_io_requestor_1_resp_bits_pte_v;
    wire ptw_io_requestor_1_resp_bits_gpa_is_pte;
    wire ptw_io_requestor_1_status_debug;
    wire ptw_io_requestor_1_pmp_0_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_0_cfg_a;
    wire ptw_io_requestor_1_pmp_0_cfg_x;
    wire ptw_io_requestor_1_pmp_0_cfg_w;
    wire ptw_io_requestor_1_pmp_0_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_0_addr;
    wire[31:0] ptw_io_requestor_1_pmp_0_mask;
    wire ptw_io_requestor_1_pmp_1_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_1_cfg_a;
    wire ptw_io_requestor_1_pmp_1_cfg_x;
    wire ptw_io_requestor_1_pmp_1_cfg_w;
    wire ptw_io_requestor_1_pmp_1_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_1_addr;
    wire[31:0] ptw_io_requestor_1_pmp_1_mask;
    wire ptw_io_requestor_1_pmp_2_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_2_cfg_a;
    wire ptw_io_requestor_1_pmp_2_cfg_x;
    wire ptw_io_requestor_1_pmp_2_cfg_w;
    wire ptw_io_requestor_1_pmp_2_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_2_addr;
    wire[31:0] ptw_io_requestor_1_pmp_2_mask;
    wire ptw_io_requestor_1_pmp_3_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_3_cfg_a;
    wire ptw_io_requestor_1_pmp_3_cfg_x;
    wire ptw_io_requestor_1_pmp_3_cfg_w;
    wire ptw_io_requestor_1_pmp_3_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_3_addr;
    wire[31:0] ptw_io_requestor_1_pmp_3_mask;
    wire ptw_io_requestor_1_pmp_4_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_4_cfg_a;
    wire ptw_io_requestor_1_pmp_4_cfg_x;
    wire ptw_io_requestor_1_pmp_4_cfg_w;
    wire ptw_io_requestor_1_pmp_4_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_4_addr;
    wire[31:0] ptw_io_requestor_1_pmp_4_mask;
    wire ptw_io_requestor_1_pmp_5_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_5_cfg_a;
    wire ptw_io_requestor_1_pmp_5_cfg_x;
    wire ptw_io_requestor_1_pmp_5_cfg_w;
    wire ptw_io_requestor_1_pmp_5_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_5_addr;
    wire[31:0] ptw_io_requestor_1_pmp_5_mask;
    wire ptw_io_requestor_1_pmp_6_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_6_cfg_a;
    wire ptw_io_requestor_1_pmp_6_cfg_x;
    wire ptw_io_requestor_1_pmp_6_cfg_w;
    wire ptw_io_requestor_1_pmp_6_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_6_addr;
    wire[31:0] ptw_io_requestor_1_pmp_6_mask;
    wire ptw_io_requestor_1_pmp_7_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_7_cfg_a;
    wire ptw_io_requestor_1_pmp_7_cfg_x;
    wire ptw_io_requestor_1_pmp_7_cfg_w;
    wire ptw_io_requestor_1_pmp_7_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_7_addr;
    wire[31:0] ptw_io_requestor_1_pmp_7_mask;
    wire[31:0] ptw_io_requestor_1_customCSRs_csrs_0_value;
    wire ptw_io_dpath_sfence_valid;
    wire ptw_io_dpath_sfence_bits_rs1;
    wire ptw_io_dpath_status_debug;
    wire ptw_io_dpath_pmp_0_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_0_cfg_a;
    wire ptw_io_dpath_pmp_0_cfg_x;
    wire ptw_io_dpath_pmp_0_cfg_w;
    wire ptw_io_dpath_pmp_0_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_0_addr;
    wire[31:0] ptw_io_dpath_pmp_0_mask;
    wire ptw_io_dpath_pmp_1_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_1_cfg_a;
    wire ptw_io_dpath_pmp_1_cfg_x;
    wire ptw_io_dpath_pmp_1_cfg_w;
    wire ptw_io_dpath_pmp_1_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_1_addr;
    wire[31:0] ptw_io_dpath_pmp_1_mask;
    wire ptw_io_dpath_pmp_2_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_2_cfg_a;
    wire ptw_io_dpath_pmp_2_cfg_x;
    wire ptw_io_dpath_pmp_2_cfg_w;
    wire ptw_io_dpath_pmp_2_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_2_addr;
    wire[31:0] ptw_io_dpath_pmp_2_mask;
    wire ptw_io_dpath_pmp_3_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_3_cfg_a;
    wire ptw_io_dpath_pmp_3_cfg_x;
    wire ptw_io_dpath_pmp_3_cfg_w;
    wire ptw_io_dpath_pmp_3_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_3_addr;
    wire[31:0] ptw_io_dpath_pmp_3_mask;
    wire ptw_io_dpath_pmp_4_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_4_cfg_a;
    wire ptw_io_dpath_pmp_4_cfg_x;
    wire ptw_io_dpath_pmp_4_cfg_w;
    wire ptw_io_dpath_pmp_4_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_4_addr;
    wire[31:0] ptw_io_dpath_pmp_4_mask;
    wire ptw_io_dpath_pmp_5_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_5_cfg_a;
    wire ptw_io_dpath_pmp_5_cfg_x;
    wire ptw_io_dpath_pmp_5_cfg_w;
    wire ptw_io_dpath_pmp_5_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_5_addr;
    wire[31:0] ptw_io_dpath_pmp_5_mask;
    wire ptw_io_dpath_pmp_6_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_6_cfg_a;
    wire ptw_io_dpath_pmp_6_cfg_x;
    wire ptw_io_dpath_pmp_6_cfg_w;
    wire ptw_io_dpath_pmp_6_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_6_addr;
    wire[31:0] ptw_io_dpath_pmp_6_mask;
    wire ptw_io_dpath_pmp_7_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_7_cfg_a;
    wire ptw_io_dpath_pmp_7_cfg_x;
    wire ptw_io_dpath_pmp_7_cfg_w;
    wire ptw_io_dpath_pmp_7_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_7_addr;
    wire[31:0] ptw_io_dpath_pmp_7_mask;
    wire[31:0] ptw_io_dpath_customCSRs_csrs_0_value;

    wire[9:0] ptw__r_pte_barrier_io_y_reserved_for_future ; 
    wire[43:0] ptw__r_pte_barrier_io_y_ppn ; 
    wire[1:0] ptw__r_pte_barrier_io_y_reserved_for_software ; 
    wire ptw__r_pte_barrier_io_y_d ; 
    wire ptw__r_pte_barrier_io_y_a ; 
    wire ptw__r_pte_barrier_io_y_g ; 
    wire ptw__r_pte_barrier_io_y_u ; 
    wire ptw__r_pte_barrier_io_y_x ; 
    wire ptw__r_pte_barrier_io_y_w ; 
    wire ptw__r_pte_barrier_io_y_r ; 
    wire ptw__r_pte_barrier_io_y_v ; 
    wire[2:0] ptw__state_barrier_io_y ; 
    wire[19:0] ptw__arb_io_out_bits_bits_addr ; 
    wire ptw__arb_io_out_bits_bits_vstage1 ; 
    wire[21:0] ptw_satp_ppn =22'h0; 
    wire[21:0] ptw_idxs_0 =22'h0; 
    wire[1:0] ptw_r_hgatp_initial_count =2'h0; 
    wire[1:0] ptw_tmp_reserved_for_software =2'h0; 
    wire[1:0] ptw_pte_reserved_for_software =2'h0; 
    wire[1:0] ptw_count_1 =2'h0; 
    wire[1:0] ptw_hits_lo_lo_1 =2'h0; 
    wire[1:0] ptw_hits_lo_hi_1 =2'h0; 
    wire[1:0] ptw_hits_hi_lo_1 =2'h0; 
    wire[1:0] ptw_hits_hi_hi_1 =2'h0; 
    wire[1:0] ptw_hi_3 =2'h0; 
    wire[1:0] ptw_lo_3 =2'h0; 
    wire[1:0] ptw_l2_pte_reserved_for_software =2'h0; 
    wire[1:0] ptw_satp_initial_count =2'h0; 
    wire[1:0] ptw_vsatp_initial_count =2'h0; 
    wire[1:0] ptw_hgatp_initial_count =2'h0; 
    wire[1:0] ptw_resp_gf_count =2'h0; 
    wire[1:0] ptw_r_pte_count =2'h0; 
    wire[1:0] ptw_r_pte_lsbs =2'h0; 
    wire[1:0] ptw_r_pte_pte_reserved_for_software =2'h0; 
    wire[1:0] ptw_r_pte_pte_1_reserved_for_software =2'h0; 
    wire[1:0] ptw_r_pte_count_1 =2'h0; 
    wire[1:0] ptw_r_pte_lsbs_1 =2'h0; 
    wire[1:0] ptw_r_pte_count_2 =2'h0; 
    wire[1:0] ptw_r_pte_idxs_0_2 =2'h0; 
    wire[1:0] ptw_r_pte_lsbs_2 =2'h0; 
    wire[1:0] ptw_aux_pte_pte_reserved_for_software =2'h0; 
    wire[3:0] ptw_hits_lo_1 =4'h0; 
    wire[3:0] ptw_hits_hi_1 =4'h0; 
    wire[3:0] ptw_hi_2 =4'h0; 
    wire[3:0] ptw_lo_2 =4'h0; 
    wire ptw_state_reg_set_left_older_9 =1'h1; 
    wire ptw_state_reg_set_left_older_10 =1'h1; 
    wire ptw_state_reg_set_left_older_11 =1'h1; 
    wire ptw_pmpHomogeneous_beginsAfterLower =1'h1; 
    wire ptw_satp_mode =1'h0; 
    wire ptw_tmp_d =1'h0; 
    wire ptw_tmp_a =1'h0; 
    wire ptw_tmp_g =1'h0; 
    wire ptw_tmp_u =1'h0; 
    wire ptw_tmp_x =1'h0; 
    wire ptw_tmp_w =1'h0; 
    wire ptw_tmp_r =1'h0; 
    wire ptw_tmp_v =1'h0; 
    wire ptw_pte_d =1'h0; 
    wire ptw_pte_a =1'h0; 
    wire ptw_pte_g =1'h0; 
    wire ptw_pte_u =1'h0; 
    wire ptw_pte_x =1'h0; 
    wire ptw_pte_w =1'h0; 
    wire ptw_pte_r =1'h0; 
    wire ptw_pte_v =1'h0; 
    wire ptw_invalid_paddr =1'h0; 
    wire ptw_invalid_gpa =1'h0; 
    wire ptw_traverse =1'h0; 
    wire ptw_stage2_pte_cache_hit =1'h0; 
    wire ptw_l2_pte_d =1'h0; 
    wire ptw_l2_pte_a =1'h0; 
    wire ptw_l2_pte_g =1'h0; 
    wire ptw_l2_pte_u =1'h0; 
    wire ptw_l2_pte_x =1'h0; 
    wire ptw_l2_pte_w =1'h0; 
    wire ptw_l2_pte_r =1'h0; 
    wire ptw_l2_pte_v =1'h0; 
    wire ptw_pmpHomogeneous_endsBeforeLower =1'h0; 
    wire ptw_do_switch =1'h0; 
    wire ptw_resp_gf_idxs_0 =1'h0; 
    wire ptw_r_pte_idxs_0 =1'h0; 
    wire ptw_r_pte_pte_d =1'h0; 
    wire ptw_r_pte_pte_a =1'h0; 
    wire ptw_r_pte_pte_g =1'h0; 
    wire ptw_r_pte_pte_u =1'h0; 
    wire ptw_r_pte_pte_x =1'h0; 
    wire ptw_r_pte_pte_w =1'h0; 
    wire ptw_r_pte_pte_r =1'h0; 
    wire ptw_r_pte_pte_v =1'h0; 
    wire ptw_r_pte_pte_1_d =1'h0; 
    wire ptw_r_pte_pte_1_a =1'h0; 
    wire ptw_r_pte_pte_1_g =1'h0; 
    wire ptw_r_pte_pte_1_u =1'h0; 
    wire ptw_r_pte_pte_1_x =1'h0; 
    wire ptw_r_pte_pte_1_w =1'h0; 
    wire ptw_r_pte_pte_1_r =1'h0; 
    wire ptw_r_pte_pte_1_v =1'h0; 
    wire ptw_ae =1'h0; 
    wire ptw_pf =1'h0; 
    wire ptw_success =1'h0; 
    wire ptw_aux_pte_pte_d =1'h0; 
    wire ptw_aux_pte_pte_a =1'h0; 
    wire ptw_aux_pte_pte_g =1'h0; 
    wire ptw_aux_pte_pte_u =1'h0; 
    wire ptw_aux_pte_pte_x =1'h0; 
    wire ptw_aux_pte_pte_w =1'h0; 
    wire ptw_aux_pte_pte_r =1'h0; 
    wire ptw_aux_pte_pte_v =1'h0; 
    wire ptw_leaf =1'h0; 
    wire ptw_leaf_1 =1'h0; 
    wire[9:0] ptw_tmp_reserved_for_future =10'h0; 
    wire[9:0] ptw_pte_reserved_for_future =10'h0; 
    wire[9:0] ptw_l2_pte_reserved_for_future =10'h0; 
    wire[9:0] ptw_r_pte_pte_reserved_for_future =10'h0; 
    wire[9:0] ptw_r_pte_pte_1_reserved_for_future =10'h0; 
    wire[9:0] ptw_aux_pte_pte_reserved_for_future =10'h0; 
    wire[43:0] ptw_tmp_ppn =44'h0; 
    wire[43:0] ptw_pte_ppn =44'h0; 
    wire[43:0] ptw_l2_pte_ppn =44'h0; 
    wire[43:0] ptw_r_pte_pte_4_ppn =44'h0; 
    wire[43:0] ptw_r_pte_pte_5_ppn =44'h0; 
    wire[8:0] ptw_satp_asid =9'h0; 
    wire[2:0] ptw_state_reg_touch_way_sized_3 =3'h0; 
    wire[23:0] ptw_r_pte_idxs_0_1 =24'h0; 
    wire[19:0] ptw_stage2_pte_cache_data =20'h0; 
    wire[7:0] ptw_hits_1 =8'h0; 
    wire[32:0] ptw_tag_1 =33'h100000000; reg[2:0] ptw_state ; 
    reg ptw_resp_valid_0 ; 
    reg ptw_resp_valid_1 ; 
    wire ptw_l2_refill_wire ; 
    wire ptw_clock_en =(| ptw_state )| ptw_l2_refill_wire | ptw_io_dpath_sfence_valid | ptw_io_dpath_customCSRs_csrs_0_value [0]; 
    reg ptw_invalidated ; 
    reg ptw_count ; 
    reg ptw_resp_ae_ptw ; 
    reg ptw_resp_ae_final ; 
    reg ptw_resp_pf ; 
    reg ptw_resp_gf ; 
    reg ptw_resp_hr ; 
    reg ptw_resp_hw ; 
    reg ptw_resp_hx ; 
    reg ptw_resp_fragmented_superpage ; reg[19:0] ptw_r_req_addr ; 
    reg ptw_r_req_need_gpa ; 
    reg ptw_r_req_vstage1 ; 
    reg ptw_r_req_stage2 ; 
    reg ptw_r_req_dest ; reg[9:0] ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_2_reserved_for_future = ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_3_reserved_for_future = ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_4_reserved_for_future = ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_5_reserved_for_future = ptw_r_pte_reserved_for_future ; reg[43:0] ptw_r_pte_ppn ; reg[1:0] ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_2_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_3_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_4_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_5_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    reg ptw_r_pte_d ; 
    wire ptw_r_pte_pte_2_d = ptw_r_pte_d ; 
    wire ptw_r_pte_pte_3_d = ptw_r_pte_d ; 
    wire ptw_r_pte_pte_4_d = ptw_r_pte_d ; 
    wire ptw_r_pte_pte_5_d = ptw_r_pte_d ; 
    reg ptw_r_pte_a ; 
    wire ptw_r_pte_pte_2_a = ptw_r_pte_a ; 
    wire ptw_r_pte_pte_3_a = ptw_r_pte_a ; 
    wire ptw_r_pte_pte_4_a = ptw_r_pte_a ; 
    wire ptw_r_pte_pte_5_a = ptw_r_pte_a ; 
    reg ptw_r_pte_g ; 
    wire ptw_r_pte_pte_2_g = ptw_r_pte_g ; 
    wire ptw_r_pte_pte_3_g = ptw_r_pte_g ; 
    wire ptw_r_pte_pte_4_g = ptw_r_pte_g ; 
    wire ptw_r_pte_pte_5_g = ptw_r_pte_g ; 
    reg ptw_r_pte_u ; 
    wire ptw_r_pte_pte_2_u = ptw_r_pte_u ; 
    wire ptw_r_pte_pte_3_u = ptw_r_pte_u ; 
    wire ptw_r_pte_pte_4_u = ptw_r_pte_u ; 
    wire ptw_r_pte_pte_5_u = ptw_r_pte_u ; 
    reg ptw_r_pte_x ; 
    wire ptw_r_pte_pte_2_x = ptw_r_pte_x ; 
    wire ptw_r_pte_pte_3_x = ptw_r_pte_x ; 
    wire ptw_r_pte_pte_4_x = ptw_r_pte_x ; 
    wire ptw_r_pte_pte_5_x = ptw_r_pte_x ; 
    reg ptw_r_pte_w ; 
    wire ptw_r_pte_pte_2_w = ptw_r_pte_w ; 
    wire ptw_r_pte_pte_3_w = ptw_r_pte_w ; 
    wire ptw_r_pte_pte_4_w = ptw_r_pte_w ; 
    wire ptw_r_pte_pte_5_w = ptw_r_pte_w ; 
    reg ptw_r_pte_r ; 
    wire ptw_r_pte_pte_2_r = ptw_r_pte_r ; 
    wire ptw_r_pte_pte_3_r = ptw_r_pte_r ; 
    wire ptw_r_pte_pte_4_r = ptw_r_pte_r ; 
    wire ptw_r_pte_pte_5_r = ptw_r_pte_r ; 
    reg ptw_r_pte_v ; 
    wire ptw_r_pte_pte_2_v = ptw_r_pte_v ; 
    wire ptw_r_pte_pte_3_v = ptw_r_pte_v ; 
    wire ptw_r_pte_pte_4_v = ptw_r_pte_v ; 
    wire ptw_r_pte_pte_5_v = ptw_r_pte_v ; 
    reg ptw_r_hgatp_mode ; reg[8:0] ptw_r_hgatp_asid ; reg[21:0] ptw_r_hgatp_ppn ; 
    reg ptw_aux_count ; reg[9:0] ptw_aux_pte_reserved_for_future ; 
    wire[9:0] ptw_merged_pte_reserved_for_future = ptw_aux_pte_reserved_for_future ; reg[43:0] ptw_aux_pte_ppn ; reg[1:0] ptw_aux_pte_reserved_for_software ; 
    wire[1:0] ptw_merged_pte_reserved_for_software = ptw_aux_pte_reserved_for_software ; 
    reg ptw_aux_pte_d ; 
    wire ptw_merged_pte_d = ptw_aux_pte_d ; 
    reg ptw_aux_pte_a ; 
    wire ptw_merged_pte_a = ptw_aux_pte_a ; 
    reg ptw_aux_pte_g ; 
    wire ptw_merged_pte_g = ptw_aux_pte_g ; 
    reg ptw_aux_pte_u ; 
    wire ptw_merged_pte_u = ptw_aux_pte_u ; 
    reg ptw_aux_pte_x ; 
    wire ptw_merged_pte_x = ptw_aux_pte_x ; 
    reg ptw_aux_pte_w ; 
    wire ptw_merged_pte_w = ptw_aux_pte_w ; 
    reg ptw_aux_pte_r ; 
    wire ptw_merged_pte_r = ptw_aux_pte_r ; 
    reg ptw_aux_pte_v ; 
    wire ptw_merged_pte_v = ptw_aux_pte_v ; reg[11:0] ptw_gpa_pgoff ; 
    reg ptw_stage2 ; 
    reg ptw_stage2_final ; 
    wire ptw_do_both_stages = ptw_r_req_vstage1 & ptw_r_req_stage2 ; 
    wire ptw_max_count = ptw_count < ptw_aux_count  ?  ptw_aux_count : ptw_count ; 
    wire[43:0] ptw_vpn = ptw_r_req_vstage1 & ptw_stage2  ?  ptw_aux_pte_ppn :{24'h0, ptw_r_req_addr }; reg[6:0] ptw_state_reg ; reg[7:0] ptw_valid ; reg[31:0] ptw_tags_0 ; reg[31:0] ptw_tags_1 ; reg[31:0] ptw_tags_2 ; reg[31:0] ptw_tags_3 ; reg[31:0] ptw_tags_4 ; reg[31:0] ptw_tags_5 ; reg[31:0] ptw_tags_6 ; reg[31:0] ptw_tags_7 ; reg[19:0] ptw_data_0 ; reg[19:0] ptw_data_1 ; reg[19:0] ptw_data_2 ; reg[19:0] ptw_data_3 ; reg[19:0] ptw_data_4 ; reg[19:0] ptw_data_5 ; reg[19:0] ptw_data_6 ; reg[19:0] ptw_data_7 ; 
    wire ptw_can_hit =~ ptw_count &( ptw_r_req_vstage1  ?  ptw_stage2 :~ ptw_r_req_stage2 ); 
    wire[32:0] ptw_tag ={ ptw_r_req_vstage1 ,32'h0}; 
    wire[1:0] ptw_hits_lo_lo ={{1'h0, ptw_tags_1 }== ptw_tag ,{1'h0, ptw_tags_0 }== ptw_tag }; 
    wire[1:0] ptw_hits_lo_hi ={{1'h0, ptw_tags_3 }== ptw_tag ,{1'h0, ptw_tags_2 }== ptw_tag }; 
    wire[3:0] ptw_hits_lo ={ ptw_hits_lo_hi , ptw_hits_lo_lo }; 
    wire[1:0] ptw_hits_hi_lo ={{1'h0, ptw_tags_5 }== ptw_tag ,{1'h0, ptw_tags_4 }== ptw_tag }; 
    wire[1:0] ptw_hits_hi_hi ={{1'h0, ptw_tags_7 }== ptw_tag ,{1'h0, ptw_tags_6 }== ptw_tag }; 
    wire[3:0] ptw_hits_hi ={ ptw_hits_hi_hi , ptw_hits_hi_lo }; 
    wire[7:0] ptw_hits ={ ptw_hits_hi , ptw_hits_lo }& ptw_valid ; 
    wire ptw_pte_cache_hit =(| ptw_hits )& ptw_can_hit ; 
    wire ptw_r_left_subtree_older = ptw_state_reg [6]; 
    wire[2:0] ptw_r_left_subtree_state = ptw_state_reg [5:3]; 
    wire[2:0] ptw_state_reg_left_subtree_state = ptw_state_reg [5:3]; 
    wire[2:0] ptw_state_reg_left_subtree_state_3 = ptw_state_reg [5:3]; 
    wire[2:0] ptw_r_right_subtree_state = ptw_state_reg [2:0]; 
    wire[2:0] ptw_state_reg_right_subtree_state = ptw_state_reg [2:0]; 
    wire[2:0] ptw_state_reg_right_subtree_state_3 = ptw_state_reg [2:0]; 
    wire ptw_r_left_subtree_older_1 = ptw_r_left_subtree_state [2]; 
    wire ptw_r_left_subtree_state_1 = ptw_r_left_subtree_state [1]; 
    wire ptw_r_right_subtree_state_1 = ptw_r_left_subtree_state [0]; 
    wire ptw_r_left_subtree_older_2 = ptw_r_right_subtree_state [2]; 
    wire ptw_r_left_subtree_state_2 = ptw_r_right_subtree_state [1]; 
    wire ptw_r_right_subtree_state_2 = ptw_r_right_subtree_state [0]; 
    wire[6:0] ptw__r_T_11 =~( ptw_valid [6:0]); 
    wire[2:0] ptw_r =(& ptw_valid ) ? { ptw_r_left_subtree_older , ptw_r_left_subtree_older  ? { ptw_r_left_subtree_older_1 , ptw_r_left_subtree_older_1  ?  ptw_r_left_subtree_state_1 : ptw_r_right_subtree_state_1 }:{ ptw_r_left_subtree_older_2 , ptw_r_left_subtree_older_2  ?  ptw_r_left_subtree_state_2 : ptw_r_right_subtree_state_2 }}: ptw__r_T_11 [0] ? 3'h0: ptw__r_T_11 [1] ? 3'h1: ptw__r_T_11 [2] ? 3'h2: ptw__r_T_11 [3] ? 3'h3: ptw__r_T_11 [4] ? 3'h4: ptw__r_T_11 [5] ? 3'h5:{2'h3,~( ptw__r_T_11 [6])}; 
    wire[2:0] ptw_state_reg_touch_way_sized = ptw_r ; 
    wire ptw_state_reg_set_left_older =~( ptw_state_reg_touch_way_sized [2]); 
    wire ptw_state_reg_set_left_older_1 =~( ptw_state_reg_touch_way_sized [1]); 
    wire ptw_state_reg_left_subtree_state_1 = ptw_state_reg_left_subtree_state [1]; 
    wire ptw_state_reg_right_subtree_state_1 = ptw_state_reg_left_subtree_state [0]; 
    wire[1:0] ptw_state_reg_hi ={ ptw_state_reg_set_left_older_1 , ptw_state_reg_set_left_older_1  ?  ptw_state_reg_left_subtree_state_1 :~( ptw_state_reg_touch_way_sized [0])}; 
    wire ptw_state_reg_set_left_older_2 =~( ptw_state_reg_touch_way_sized [1]); 
    wire ptw_state_reg_left_subtree_state_2 = ptw_state_reg_right_subtree_state [1]; 
    wire ptw_state_reg_right_subtree_state_2 = ptw_state_reg_right_subtree_state [0]; 
    wire[1:0] ptw_state_reg_hi_1 ={ ptw_state_reg_set_left_older_2 , ptw_state_reg_set_left_older_2  ?  ptw_state_reg_left_subtree_state_2 :~( ptw_state_reg_touch_way_sized [0])}; 
    wire[3:0] ptw_state_reg_hi_2 ={ ptw_state_reg_set_left_older , ptw_state_reg_set_left_older  ?  ptw_state_reg_left_subtree_state :{ ptw_state_reg_hi , ptw_state_reg_set_left_older_1  ? ~( ptw_state_reg_touch_way_sized [0]): ptw_state_reg_right_subtree_state_1 }}; 
    wire ptw__r_pte_T_6 = ptw_state ==3'h1; 
    wire[3:0] ptw_hi = ptw_hits [7:4]; 
    wire[3:0] ptw_lo = ptw_hits [3:0]; 
    wire[3:0] ptw__GEN = ptw_hi | ptw_lo ; 
    wire[1:0] ptw_hi_1 = ptw__GEN [3:2]; 
    wire[1:0] ptw_lo_1 = ptw__GEN [1:0]; 
    wire[2:0] ptw_state_reg_touch_way_sized_1 ={| ptw_hi ,| ptw_hi_1 , ptw_hi_1 [1]| ptw_lo_1 [1]}; 
    wire ptw_state_reg_set_left_older_3 =~( ptw_state_reg_touch_way_sized_1 [2]); 
    wire ptw_state_reg_set_left_older_4 =~( ptw_state_reg_touch_way_sized_1 [1]); 
    wire ptw_state_reg_left_subtree_state_4 = ptw_state_reg_left_subtree_state_3 [1]; 
    wire ptw_state_reg_right_subtree_state_4 = ptw_state_reg_left_subtree_state_3 [0]; 
    wire[1:0] ptw_state_reg_hi_3 ={ ptw_state_reg_set_left_older_4 , ptw_state_reg_set_left_older_4  ?  ptw_state_reg_left_subtree_state_4 :~( ptw_state_reg_touch_way_sized_1 [0])}; 
    wire ptw_state_reg_set_left_older_5 =~( ptw_state_reg_touch_way_sized_1 [1]); 
    wire ptw_state_reg_left_subtree_state_5 = ptw_state_reg_right_subtree_state_3 [1]; 
    wire ptw_state_reg_right_subtree_state_5 = ptw_state_reg_right_subtree_state_3 [0]; 
    wire[1:0] ptw_state_reg_hi_4 ={ ptw_state_reg_set_left_older_5 , ptw_state_reg_set_left_older_5  ?  ptw_state_reg_left_subtree_state_5 :~( ptw_state_reg_touch_way_sized_1 [0])}; 
    wire[3:0] ptw_state_reg_hi_5 ={ ptw_state_reg_set_left_older_3 , ptw_state_reg_set_left_older_3  ?  ptw_state_reg_left_subtree_state_3 :{ ptw_state_reg_hi_3 , ptw_state_reg_set_left_older_4  ? ~( ptw_state_reg_touch_way_sized_1 [0]): ptw_state_reg_right_subtree_state_4 }}; 
    wire[19:0] ptw_pte_cache_data =( ptw_hits [0] ?  ptw_data_0 :20'h0)|( ptw_hits [1] ?  ptw_data_1 :20'h0)|( ptw_hits [2] ?  ptw_data_2 :20'h0)|( ptw_hits [3] ?  ptw_data_3 :20'h0)|( ptw_hits [4] ?  ptw_data_4 :20'h0)|( ptw_hits [5] ?  ptw_data_5 :20'h0)|( ptw_hits [6] ?  ptw_data_6 :20'h0)|( ptw_hits [7] ?  ptw_data_7 :20'h0); reg[6:0] ptw_state_reg_1 ; reg[7:0] ptw_valid_1 ; reg[19:0] ptw_data_1_0 ; reg[19:0] ptw_data_1_1 ; reg[19:0] ptw_data_1_2 ; reg[19:0] ptw_data_1_3 ; reg[19:0] ptw_data_1_4 ; reg[19:0] ptw_data_1_5 ; reg[19:0] ptw_data_1_6 ; reg[19:0] ptw_data_1_7 ; 
    wire ptw_can_hit_1 =~ ptw_count &~ ptw_aux_count & ptw_r_req_vstage1 & ptw_stage2 &~ ptw_stage2_final ; 
    wire ptw_can_refill = ptw_do_both_stages &~ ptw_stage2 &~ ptw_stage2_final ; 
    wire ptw_r_left_subtree_older_3 = ptw_state_reg_1 [6]; 
    wire[2:0] ptw_r_left_subtree_state_3 = ptw_state_reg_1 [5:3]; 
    wire[2:0] ptw_state_reg_left_subtree_state_6 = ptw_state_reg_1 [5:3]; 
    wire[2:0] ptw_state_reg_left_subtree_state_9 = ptw_state_reg_1 [5:3]; 
    wire[2:0] ptw_r_right_subtree_state_3 = ptw_state_reg_1 [2:0]; 
    wire[2:0] ptw_state_reg_right_subtree_state_6 = ptw_state_reg_1 [2:0]; 
    wire[2:0] ptw_state_reg_right_subtree_state_9 = ptw_state_reg_1 [2:0]; 
    wire ptw_r_left_subtree_older_4 = ptw_r_left_subtree_state_3 [2]; 
    wire ptw_r_left_subtree_state_4 = ptw_r_left_subtree_state_3 [1]; 
    wire ptw_r_right_subtree_state_4 = ptw_r_left_subtree_state_3 [0]; 
    wire ptw_r_left_subtree_older_5 = ptw_r_right_subtree_state_3 [2]; 
    wire ptw_r_left_subtree_state_5 = ptw_r_right_subtree_state_3 [1]; 
    wire ptw_r_right_subtree_state_5 = ptw_r_right_subtree_state_3 [0]; 
    wire[6:0] ptw__r_T_38 =~( ptw_valid_1 [6:0]); 
    wire[2:0] ptw_r_1 =(& ptw_valid_1 ) ? { ptw_r_left_subtree_older_3 , ptw_r_left_subtree_older_3  ? { ptw_r_left_subtree_older_4 , ptw_r_left_subtree_older_4  ?  ptw_r_left_subtree_state_4 : ptw_r_right_subtree_state_4 }:{ ptw_r_left_subtree_older_5 , ptw_r_left_subtree_older_5  ?  ptw_r_left_subtree_state_5 : ptw_r_right_subtree_state_5 }}: ptw__r_T_38 [0] ? 3'h0: ptw__r_T_38 [1] ? 3'h1: ptw__r_T_38 [2] ? 3'h2: ptw__r_T_38 [3] ? 3'h3: ptw__r_T_38 [4] ? 3'h4: ptw__r_T_38 [5] ? 3'h5:{2'h3,~( ptw__r_T_38 [6])}; 
    wire[2:0] ptw_state_reg_touch_way_sized_2 = ptw_r_1 ; 
    wire ptw_state_reg_set_left_older_6 =~( ptw_state_reg_touch_way_sized_2 [2]); 
    wire ptw_state_reg_set_left_older_7 =~( ptw_state_reg_touch_way_sized_2 [1]); 
    wire ptw_state_reg_left_subtree_state_7 = ptw_state_reg_left_subtree_state_6 [1]; 
    wire ptw_state_reg_right_subtree_state_7 = ptw_state_reg_left_subtree_state_6 [0]; 
    wire[1:0] ptw_state_reg_hi_6 ={ ptw_state_reg_set_left_older_7 , ptw_state_reg_set_left_older_7  ?  ptw_state_reg_left_subtree_state_7 :~( ptw_state_reg_touch_way_sized_2 [0])}; 
    wire ptw_state_reg_set_left_older_8 =~( ptw_state_reg_touch_way_sized_2 [1]); 
    wire ptw_state_reg_left_subtree_state_8 = ptw_state_reg_right_subtree_state_6 [1]; 
    wire ptw_state_reg_right_subtree_state_8 = ptw_state_reg_right_subtree_state_6 [0]; 
    wire[1:0] ptw_state_reg_hi_7 ={ ptw_state_reg_set_left_older_8 , ptw_state_reg_set_left_older_8  ?  ptw_state_reg_left_subtree_state_8 :~( ptw_state_reg_touch_way_sized_2 [0])}; 
    wire[3:0] ptw_state_reg_hi_8 ={ ptw_state_reg_set_left_older_6 , ptw_state_reg_set_left_older_6  ?  ptw_state_reg_left_subtree_state_6 :{ ptw_state_reg_hi_6 , ptw_state_reg_set_left_older_7  ? ~( ptw_state_reg_touch_way_sized_2 [0]): ptw_state_reg_right_subtree_state_7 }}; 
    wire ptw_state_reg_left_subtree_state_10 = ptw_state_reg_left_subtree_state_9 [1]; 
    wire ptw_state_reg_right_subtree_state_10 = ptw_state_reg_left_subtree_state_9 [0]; 
    wire[1:0] ptw_state_reg_hi_9 ={1'h1, ptw_state_reg_left_subtree_state_10 }; 
    wire ptw_state_reg_left_subtree_state_11 = ptw_state_reg_right_subtree_state_9 [1]; 
    wire ptw_state_reg_right_subtree_state_11 = ptw_state_reg_right_subtree_state_9 [0]; 
    wire[1:0] ptw_state_reg_hi_10 ={1'h1, ptw_state_reg_left_subtree_state_11 }; 
    wire[3:0] ptw_state_reg_hi_11 ={1'h1, ptw_state_reg_left_subtree_state_9 }; 
    reg ptw_pte_hit ; 
    reg ptw_l2_refill ; 
  assign  ptw_l2_refill_wire = ptw_l2_refill ; 
    wire[55:0] ptw__pmpHomogeneous_T ={ ptw_r_pte_ppn ,12'h0}; 
    wire[29:0] ptw__GEN_0 ={ ptw_r_pte_ppn [43:16],~( ptw_r_pte_ppn [15:14])}; 
    wire[26:0] ptw__GEN_1 ={ ptw_r_pte_ppn [43:19],~( ptw_r_pte_ppn [18:17])}; 
    wire ptw_pmaPgLevelHomogeneous_0 = ptw__GEN_0 ==30'h0| ptw__GEN_1 ==27'h0; 
    wire[31:0] ptw__GEN_2 ={ ptw_r_pte_ppn [19:0],12'h0}; 
    wire ptw_pmaPgLevelHomogeneous_1 = ptw_r_pte_ppn ==44'h0|{ ptw_r_pte_ppn [43:2],~( ptw_r_pte_ppn [1:0])}==44'h0|{ ptw_r_pte_ppn [43:5],~( ptw_r_pte_ppn [4])}==40'h0|{ ptw_r_pte_ppn [43:14], ptw_r_pte_ppn [13:4]^10'h200}==40'h0| ptw__GEN_0 ==30'h0| ptw__GEN_1 ==27'h0|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:2]^18'h20000}==42'h0; 
    wire ptw_pmaHomogeneous = ptw_count  ?  ptw_pmaPgLevelHomogeneous_1 : ptw_pmaPgLevelHomogeneous_0 ; 
    wire ptw_pmpHomogeneous_maskHomogeneous = ptw_count  ?  ptw_io_dpath_pmp_0_mask [11]: ptw_io_dpath_pmp_0_mask [21]; 
    wire ptw__GEN_3 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_0_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper = ptw__GEN_3 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_1 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_1 = ptw__GEN_3 ; 
    wire[31:0] ptw__GEN_4 = ptw_count  ? 32'hFFFFF000:32'hFFC00000; 
    wire[31:0] ptw_pmpHomogeneous_pgMask ; 
  assign  ptw_pmpHomogeneous_pgMask = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_1 ; 
  assign  ptw_pmpHomogeneous_pgMask_1 = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_2 ; 
  assign  ptw_pmpHomogeneous_pgMask_2 = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_3 ; 
  assign  ptw_pmpHomogeneous_pgMask_3 = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_4 ; 
  assign  ptw_pmpHomogeneous_pgMask_4 = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_5 ; 
  assign  ptw_pmpHomogeneous_pgMask_5 = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_6 ; 
  assign  ptw_pmpHomogeneous_pgMask_6 = ptw__GEN_4 ; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_7 ; 
  assign  ptw_pmpHomogeneous_pgMask_7 = ptw__GEN_4 ; 
    wire ptw_pmpHomogeneous_endsBeforeUpper =( ptw__GEN_2 & ptw_pmpHomogeneous_pgMask )<({ ptw_io_dpath_pmp_0_addr ,2'h0}& ptw_pmpHomogeneous_pgMask ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_1 = ptw_count  ?  ptw_io_dpath_pmp_1_mask [11]: ptw_io_dpath_pmp_1_mask [21]; 
    wire ptw__GEN_5 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_1_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_1 ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper_1 = ptw__GEN_5 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_2 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_2 = ptw__GEN_5 ; 
    wire[31:0] ptw__GEN_6 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_1 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_1 = ptw__GEN_6 <({ ptw_io_dpath_pmp_0_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_1 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_1 = ptw__GEN_6 <({ ptw_io_dpath_pmp_1_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_1 ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_2 = ptw_count  ?  ptw_io_dpath_pmp_2_mask [11]: ptw_io_dpath_pmp_2_mask [21]; 
    wire ptw__GEN_7 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_2_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_2 ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper_2 = ptw__GEN_7 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_3 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_3 = ptw__GEN_7 ; 
    wire[31:0] ptw__GEN_8 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_2 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_2 = ptw__GEN_8 <({ ptw_io_dpath_pmp_1_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_2 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_2 = ptw__GEN_8 <({ ptw_io_dpath_pmp_2_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_2 ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_3 = ptw_count  ?  ptw_io_dpath_pmp_3_mask [11]: ptw_io_dpath_pmp_3_mask [21]; 
    wire ptw__GEN_9 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_3_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_3 ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper_3 = ptw__GEN_9 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_4 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_4 = ptw__GEN_9 ; 
    wire[31:0] ptw__GEN_10 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_3 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_3 = ptw__GEN_10 <({ ptw_io_dpath_pmp_2_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_3 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_3 = ptw__GEN_10 <({ ptw_io_dpath_pmp_3_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_3 ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_4 = ptw_count  ?  ptw_io_dpath_pmp_4_mask [11]: ptw_io_dpath_pmp_4_mask [21]; 
    wire ptw__GEN_11 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_4_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_4 ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper_4 = ptw__GEN_11 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_5 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_5 = ptw__GEN_11 ; 
    wire[31:0] ptw__GEN_12 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_4 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_4 = ptw__GEN_12 <({ ptw_io_dpath_pmp_3_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_4 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_4 = ptw__GEN_12 <({ ptw_io_dpath_pmp_4_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_4 ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_5 = ptw_count  ?  ptw_io_dpath_pmp_5_mask [11]: ptw_io_dpath_pmp_5_mask [21]; 
    wire ptw__GEN_13 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_5_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_5 ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper_5 = ptw__GEN_13 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_6 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_6 = ptw__GEN_13 ; 
    wire[31:0] ptw__GEN_14 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_5 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_5 = ptw__GEN_14 <({ ptw_io_dpath_pmp_4_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_5 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_5 = ptw__GEN_14 <({ ptw_io_dpath_pmp_5_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_5 ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_6 = ptw_count  ?  ptw_io_dpath_pmp_6_mask [11]: ptw_io_dpath_pmp_6_mask [21]; 
    wire ptw__GEN_15 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_6_addr ,2'h0}; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_6 ; 
  assign  ptw_pmpHomogeneous_beginsAfterUpper_6 = ptw__GEN_15 ; 
    wire ptw_pmpHomogeneous_beginsAfterLower_7 ; 
  assign  ptw_pmpHomogeneous_beginsAfterLower_7 = ptw__GEN_15 ; 
    wire[31:0] ptw__GEN_16 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_6 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_6 = ptw__GEN_16 <({ ptw_io_dpath_pmp_5_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_6 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_6 = ptw__GEN_16 <({ ptw_io_dpath_pmp_6_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_6 ); 
    wire ptw_pmpHomogeneous_maskHomogeneous_7 = ptw_count  ?  ptw_io_dpath_pmp_7_mask [11]: ptw_io_dpath_pmp_7_mask [21]; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_7 = ptw__pmpHomogeneous_T >={24'h0, ptw_io_dpath_pmp_7_addr ,2'h0}; 
    wire[31:0] ptw__GEN_17 = ptw__GEN_2 & ptw_pmpHomogeneous_pgMask_7 ; 
    wire ptw_pmpHomogeneous_endsBeforeLower_7 = ptw__GEN_17 <({ ptw_io_dpath_pmp_6_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_7 ); 
    wire ptw_pmpHomogeneous_endsBeforeUpper_7 = ptw__GEN_17 <({ ptw_io_dpath_pmp_7_addr ,2'h0}& ptw_pmpHomogeneous_pgMask_7 ); 
    wire ptw_pmpHomogeneous =( ptw_io_dpath_pmp_0_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_0_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_0_addr [29:20]})):~( ptw_io_dpath_pmp_0_cfg_a [0])| ptw_pmpHomogeneous_beginsAfterUpper | ptw_pmpHomogeneous_endsBeforeUpper )&( ptw_io_dpath_pmp_1_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_1 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_1_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_1_addr [29:20]})):~( ptw_io_dpath_pmp_1_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_1 | ptw_pmpHomogeneous_beginsAfterUpper_1 | ptw_pmpHomogeneous_beginsAfterLower_1 & ptw_pmpHomogeneous_endsBeforeUpper_1 )&( ptw_io_dpath_pmp_2_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_2 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_2_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_2_addr [29:20]})):~( ptw_io_dpath_pmp_2_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_2 | ptw_pmpHomogeneous_beginsAfterUpper_2 | ptw_pmpHomogeneous_beginsAfterLower_2 & ptw_pmpHomogeneous_endsBeforeUpper_2 )&( ptw_io_dpath_pmp_3_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_3 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_3_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_3_addr [29:20]})):~( ptw_io_dpath_pmp_3_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_3 | ptw_pmpHomogeneous_beginsAfterUpper_3 | ptw_pmpHomogeneous_beginsAfterLower_3 & ptw_pmpHomogeneous_endsBeforeUpper_3 )&( ptw_io_dpath_pmp_4_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_4 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_4_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_4_addr [29:20]})):~( ptw_io_dpath_pmp_4_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_4 | ptw_pmpHomogeneous_beginsAfterUpper_4 | ptw_pmpHomogeneous_beginsAfterLower_4 & ptw_pmpHomogeneous_endsBeforeUpper_4 )&( ptw_io_dpath_pmp_5_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_5 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_5_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_5_addr [29:20]})):~( ptw_io_dpath_pmp_5_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_5 | ptw_pmpHomogeneous_beginsAfterUpper_5 | ptw_pmpHomogeneous_beginsAfterLower_5 & ptw_pmpHomogeneous_endsBeforeUpper_5 )&( ptw_io_dpath_pmp_6_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_6 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_6_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_6_addr [29:20]})):~( ptw_io_dpath_pmp_6_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_6 | ptw_pmpHomogeneous_beginsAfterUpper_6 | ptw_pmpHomogeneous_beginsAfterLower_6 & ptw_pmpHomogeneous_endsBeforeUpper_6 )&( ptw_io_dpath_pmp_7_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_7 |( ptw_count  ? (|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:0]^ ptw_io_dpath_pmp_7_addr [29:10]}):(|{ ptw_r_pte_ppn [43:20], ptw_r_pte_ppn [19:10]^ ptw_io_dpath_pmp_7_addr [29:20]})):~( ptw_io_dpath_pmp_7_cfg_a [0])| ptw_pmpHomogeneous_endsBeforeLower_7 | ptw_pmpHomogeneous_beginsAfterUpper_7 | ptw_pmpHomogeneous_beginsAfterLower_7 & ptw_pmpHomogeneous_endsBeforeUpper_7 ); 
    wire ptw_homogeneous = ptw_pmaHomogeneous & ptw_pmpHomogeneous ; 
    wire[21:0] ptw_aux_ppn = ptw__arb_io_out_bits_bits_vstage1  ? 22'h0:{2'h0, ptw__arb_io_out_bits_bits_addr }; reg[2:0] ptw_casez_tmp ; 
  always @(*)
         begin 
             casez ( ptw_state )
              3 'b000: 
                  ptw_casez_tmp  = ptw_state ;
              3 'b001: 
                  ptw_casez_tmp  = ptw_resp_gf  ? 3'h0: ptw_pte_cache_hit  ?  ptw_state :3'h1;
              3 'b010: 
                  ptw_casez_tmp  =3'h4;
              3 'b011: 
                  ptw_casez_tmp  = ptw_state ;
              3 'b100: 
                  ptw_casez_tmp  =3'h5;
              3 'b101: 
                  ptw_casez_tmp  = ptw_state ;
              3 'b110: 
                  ptw_casez_tmp  = ptw_state ;
              default : 
                  ptw_casez_tmp  =3'h0;endcase
         end
    wire[2:0] ptw_next_state = ptw_casez_tmp ; 
    wire[43:0] ptw_merged_pte_superpage_mask =~ ptw_stage2_final | ptw_max_count  ? 44'hFFFFFFFFFFF:44'hFFFFFFFFC00; 
    wire[43:0] ptw_merged_pte_stage1_ppns_0 ={34'h0, ptw_aux_pte_ppn [9:0]}; 
    wire[43:0] ptw_merged_pte_stage1_ppn = ptw_count  ? 44'h0: ptw_merged_pte_stage1_ppns_0 ; 
    wire[43:0] ptw_merged_pte_ppn = ptw_merged_pte_stage1_ppn & ptw_merged_pte_superpage_mask ; 
    wire[43:0] ptw__GEN_18 ={22'h0, ptw_r_hgatp_ppn [21:2],2'h0}; 
    wire[43:0] ptw_r_pte_pte_ppn ; 
  assign  ptw_r_pte_pte_ppn = ptw__GEN_18 ; 
    wire[43:0] ptw_r_pte_pte_2_ppn ; 
  assign  ptw_r_pte_pte_2_ppn = ptw__GEN_18 ; 
    wire ptw__r_pte_T_7 = ptw__r_pte_T_6 & ptw_pte_cache_hit ; 
    wire[43:0] ptw_r_pte_pte_1_ppn ={24'h0, ptw_pte_cache_data }; 
    wire ptw__r_pte_T_16 =(& ptw_state )&~ ptw_homogeneous &~ ptw_count ; 
    wire[43:0] ptw_r_pte_pte_3_ppn ={ ptw_r_pte_ppn [43:10], ptw_r_req_addr [9:0]}; 
    wire ptw_gf = ptw_stage2 &~ ptw_stage2_final ; 
    wire[43:0] ptw_aux_pte_s1_ppns_0 ={34'h0, ptw_r_req_addr [9:0]}; 
    wire[43:0] ptw_aux_pte_pte_ppn = ptw_count  ? 44'h0: ptw_aux_pte_s1_ppns_0 ; 
    wire ptw__GEN_19 = ptw_state ==3'h0; 
    wire ptw__GEN_20 = ptw_state ==3'h1; 
    wire ptw__GEN_21 = ptw_state ==3'h2| ptw_state ==3'h4; 
  always @( posedge  ptw_clock )
         begin 
             if ( ptw_reset )
                 begin  
                     ptw_state  <=3'h0; 
                     ptw_state_reg  <=7'h0; 
                     ptw_valid  <=8'h0; 
                     ptw_state_reg_1  <=7'h0; 
                     ptw_valid_1  <=8'h0;
                 end 
              else 
                 begin  
                     ptw_state  <= ptw__state_barrier_io_y ;
                     if ( ptw_pte_cache_hit & ptw__r_pte_T_6 ) 
                         ptw_state_reg  <={ ptw_state_reg_hi_5 , ptw_state_reg_set_left_older_3  ? { ptw_state_reg_hi_4 , ptw_state_reg_set_left_older_5  ? ~( ptw_state_reg_touch_way_sized_1 [0]): ptw_state_reg_right_subtree_state_5 }: ptw_state_reg_right_subtree_state_3 };
                     if ( ptw_io_dpath_sfence_valid &~ ptw_io_dpath_sfence_bits_rs1 )
                         begin  
                             ptw_valid  <=8'h0; 
                             ptw_valid_1  <=8'h0;
                         end 
                 end  
             ptw_resp_valid_0  <=~ ptw__GEN_19 &( ptw__GEN_20  ?  ptw_resp_gf &~ ptw_r_req_dest :~ ptw__GEN_21 &(& ptw_state )&~ ptw_r_req_dest ); 
             ptw_resp_valid_1  <=~ ptw__GEN_19 &( ptw__GEN_20  ?  ptw_resp_gf & ptw_r_req_dest :~ ptw__GEN_21 &(& ptw_state )& ptw_r_req_dest ); 
             ptw_invalidated  <= ptw_io_dpath_sfence_valid | ptw_invalidated &(| ptw_state );
             if (~ ptw__GEN_19 )
                 begin 
                     if ( ptw__GEN_20 )
                         begin 
                             if ( ptw_pte_cache_hit ) 
                                 ptw_count  <= ptw_count -1'h1;
                         end 
                      else  
                         ptw_count  <=~ ptw__GEN_21 &(& ptw_state )&~ ptw_homogeneous | ptw_count ;
                 end  
             ptw_resp_fragmented_superpage  <=~ ptw__GEN_19 &~( ptw__GEN_20 | ptw__GEN_21 )&(& ptw_state )&( ptw_do_both_stages |~ ptw_homogeneous )| ptw_resp_fragmented_superpage ; 
             ptw_r_pte_reserved_for_future  <= ptw__r_pte_barrier_io_y_reserved_for_future ; 
             ptw_r_pte_ppn  <= ptw__r_pte_barrier_io_y_ppn ; 
             ptw_r_pte_reserved_for_software  <= ptw__r_pte_barrier_io_y_reserved_for_software ; 
             ptw_r_pte_d  <= ptw__r_pte_barrier_io_y_d ; 
             ptw_r_pte_a  <= ptw__r_pte_barrier_io_y_a ; 
             ptw_r_pte_g  <= ptw__r_pte_barrier_io_y_g ; 
             ptw_r_pte_u  <= ptw__r_pte_barrier_io_y_u ; 
             ptw_r_pte_x  <= ptw__r_pte_barrier_io_y_x ; 
             ptw_r_pte_w  <= ptw__r_pte_barrier_io_y_w ; 
             ptw_r_pte_r  <= ptw__r_pte_barrier_io_y_r ; 
             ptw_r_pte_v  <= ptw__r_pte_barrier_io_y_v ;
             if ( ptw__GEN_19 |~( ptw__GEN_20 & ptw_stage2 &~ ptw_count ))
                 begin 
                 end 
              else  
                 ptw_gpa_pgoff  <= ptw_aux_count  ? { ptw_r_req_addr [9:0],2'h0}:12'h0; 
             ptw_pte_hit  <=~ ptw__GEN_19 & ptw__GEN_20 & ptw_pte_cache_hit ; 
             ptw_l2_refill  <=1'h0;
         end
    wire[19:0] ptw_arb_io_in_0_bits_bits_addr;
    wire ptw_arb_io_in_0_bits_bits_need_gpa;
    wire ptw_arb_io_in_0_bits_bits_vstage1;
    wire ptw_arb_io_in_0_bits_bits_stage2;
    wire ptw_arb_io_in_1_bits_valid;
    wire[19:0] ptw_arb_io_in_1_bits_bits_addr;
    wire ptw_arb_io_in_1_bits_bits_need_gpa;
    wire ptw_arb_io_in_1_bits_bits_vstage1;
    wire ptw_arb_io_in_1_bits_bits_stage2;
    wire ptw_arb_io_out_bits_valid;
    wire[19:0] ptw_arb_io_out_bits_bits_addr;
    wire ptw_arb_io_out_bits_bits_need_gpa;
    wire ptw_arb_io_out_bits_bits_vstage1;
    wire ptw_arb_io_out_bits_bits_stage2;

    wire ptw_arb_grant_1 =1'h1; 
  assign  ptw_arb_io_out_bits_valid = ptw_arb_io_in_1_bits_valid ; 
  assign  ptw_arb_io_out_bits_bits_addr = ptw_arb_io_in_1_bits_bits_addr ; 
  assign  ptw_arb_io_out_bits_bits_need_gpa = ptw_arb_io_in_1_bits_bits_need_gpa ; 
  assign  ptw_arb_io_out_bits_bits_vstage1 = ptw_arb_io_in_1_bits_bits_vstage1 ; 
  assign  ptw_arb_io_out_bits_bits_stage2 = ptw_arb_io_in_1_bits_bits_stage2 ;
    assign ptw_arb_io_in_0_bits_bits_addr = ptw_io_requestor_0_req_bits_bits_addr;
    assign ptw_arb_io_in_0_bits_bits_need_gpa = ptw_io_requestor_0_req_bits_bits_need_gpa;
    assign ptw_arb_io_in_0_bits_bits_vstage1 = ptw_io_requestor_0_req_bits_bits_vstage1;
    assign ptw_arb_io_in_0_bits_bits_stage2 = ptw_io_requestor_0_req_bits_bits_stage2;
    assign ptw_arb_io_in_1_bits_valid = ptw_io_requestor_1_req_bits_valid;
    assign ptw_arb_io_in_1_bits_bits_addr = ptw_io_requestor_1_req_bits_bits_addr;
    assign ptw_arb_io_in_1_bits_bits_need_gpa = ptw_io_requestor_1_req_bits_bits_need_gpa;
    assign ptw_arb_io_in_1_bits_bits_vstage1 = ptw_io_requestor_1_req_bits_bits_vstage1;
    assign ptw_arb_io_in_1_bits_bits_stage2 = ptw_io_requestor_1_req_bits_bits_stage2;
    assign ptw__arb_io_out_bits_bits_addr = ptw_arb_io_out_bits_bits_addr;
    assign ptw__arb_io_out_bits_bits_vstage1 = ptw_arb_io_out_bits_bits_vstage1;
      
    wire[2:0] ptw_state_barrier_io_x;
    wire[2:0] ptw_state_barrier_io_y;

    assign  ptw_state_barrier_io_y = ptw_state_barrier_io_x ;
    assign ptw_state_barrier_io_x = ptw_next_state;
    assign ptw__state_barrier_io_y = ptw_state_barrier_io_y;
      
    wire[9:0] ptw_r_pte_barrier_io_x_reserved_for_future;
    wire[43:0] ptw_r_pte_barrier_io_x_ppn;
    wire[1:0] ptw_r_pte_barrier_io_x_reserved_for_software;
    wire ptw_r_pte_barrier_io_x_d;
    wire ptw_r_pte_barrier_io_x_a;
    wire ptw_r_pte_barrier_io_x_g;
    wire ptw_r_pte_barrier_io_x_u;
    wire ptw_r_pte_barrier_io_x_x;
    wire ptw_r_pte_barrier_io_x_w;
    wire ptw_r_pte_barrier_io_x_r;
    wire ptw_r_pte_barrier_io_x_v;
    wire[9:0] ptw_r_pte_barrier_io_y_reserved_for_future;
    wire[43:0] ptw_r_pte_barrier_io_y_ppn;
    wire[1:0] ptw_r_pte_barrier_io_y_reserved_for_software;
    wire ptw_r_pte_barrier_io_y_d;
    wire ptw_r_pte_barrier_io_y_a;
    wire ptw_r_pte_barrier_io_y_g;
    wire ptw_r_pte_barrier_io_y_u;
    wire ptw_r_pte_barrier_io_y_x;
    wire ptw_r_pte_barrier_io_y_w;
    wire ptw_r_pte_barrier_io_y_r;
    wire ptw_r_pte_barrier_io_y_v;

    assign  ptw_r_pte_barrier_io_y_reserved_for_future = ptw_r_pte_barrier_io_x_reserved_for_future ; 
  assign  ptw_r_pte_barrier_io_y_ppn = ptw_r_pte_barrier_io_x_ppn ; 
  assign  ptw_r_pte_barrier_io_y_reserved_for_software = ptw_r_pte_barrier_io_x_reserved_for_software ; 
  assign  ptw_r_pte_barrier_io_y_d = ptw_r_pte_barrier_io_x_d ; 
  assign  ptw_r_pte_barrier_io_y_a = ptw_r_pte_barrier_io_x_a ; 
  assign  ptw_r_pte_barrier_io_y_g = ptw_r_pte_barrier_io_x_g ; 
  assign  ptw_r_pte_barrier_io_y_u = ptw_r_pte_barrier_io_x_u ; 
  assign  ptw_r_pte_barrier_io_y_x = ptw_r_pte_barrier_io_x_x ; 
  assign  ptw_r_pte_barrier_io_y_w = ptw_r_pte_barrier_io_x_w ; 
  assign  ptw_r_pte_barrier_io_y_r = ptw_r_pte_barrier_io_x_r ; 
  assign  ptw_r_pte_barrier_io_y_v = ptw_r_pte_barrier_io_x_v ;
    assign ptw_r_pte_barrier_io_x_reserved_for_future = ptw__r_pte_T_7 ? 10'h0:ptw__r_pte_T_16 ? ptw_r_pte_pte_3_reserved_for_future:ptw_r_pte_reserved_for_future;
    assign ptw_r_pte_barrier_io_x_ppn = ptw__r_pte_T_7 ? ptw_r_pte_pte_1_ppn:ptw__r_pte_T_16 ? ptw_r_pte_pte_3_ppn:ptw_r_pte_ppn;
    assign ptw_r_pte_barrier_io_x_reserved_for_software = ptw__r_pte_T_7 ? 2'h0:ptw__r_pte_T_16 ? ptw_r_pte_pte_3_reserved_for_software:ptw_r_pte_reserved_for_software;
    assign ptw_r_pte_barrier_io_x_d = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_d:ptw_r_pte_d);
    assign ptw_r_pte_barrier_io_x_a = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_a:ptw_r_pte_a);
    assign ptw_r_pte_barrier_io_x_g = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_g:ptw_r_pte_g);
    assign ptw_r_pte_barrier_io_x_u = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_u:ptw_r_pte_u);
    assign ptw_r_pte_barrier_io_x_x = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_x:ptw_r_pte_x);
    assign ptw_r_pte_barrier_io_x_w = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_w:ptw_r_pte_w);
    assign ptw_r_pte_barrier_io_x_r = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_r:ptw_r_pte_r);
    assign ptw_r_pte_barrier_io_x_v = ~ptw__r_pte_T_7&(ptw__r_pte_T_16 ? ptw_r_pte_pte_3_v:ptw_r_pte_v);
    assign ptw__r_pte_barrier_io_y_reserved_for_future = ptw_r_pte_barrier_io_y_reserved_for_future;
    assign ptw__r_pte_barrier_io_y_ppn = ptw_r_pte_barrier_io_y_ppn;
    assign ptw__r_pte_barrier_io_y_reserved_for_software = ptw_r_pte_barrier_io_y_reserved_for_software;
    assign ptw__r_pte_barrier_io_y_d = ptw_r_pte_barrier_io_y_d;
    assign ptw__r_pte_barrier_io_y_a = ptw_r_pte_barrier_io_y_a;
    assign ptw__r_pte_barrier_io_y_g = ptw_r_pte_barrier_io_y_g;
    assign ptw__r_pte_barrier_io_y_u = ptw_r_pte_barrier_io_y_u;
    assign ptw__r_pte_barrier_io_y_x = ptw_r_pte_barrier_io_y_x;
    assign ptw__r_pte_barrier_io_y_w = ptw_r_pte_barrier_io_y_w;
    assign ptw__r_pte_barrier_io_y_r = ptw_r_pte_barrier_io_y_r;
    assign ptw__r_pte_barrier_io_y_v = ptw_r_pte_barrier_io_y_v;
     
  assign  ptw_io_requestor_0_resp_bits_ae_ptw = ptw_resp_ae_ptw ; 
  assign  ptw_io_requestor_0_resp_bits_ae_final = ptw_resp_ae_final ; 
  assign  ptw_io_requestor_0_resp_bits_pf = ptw_resp_pf ; 
  assign  ptw_io_requestor_0_resp_bits_gf = ptw_resp_gf ; 
  assign  ptw_io_requestor_0_resp_bits_hr = ptw_resp_hr ; 
  assign  ptw_io_requestor_0_resp_bits_hw = ptw_resp_hw ; 
  assign  ptw_io_requestor_0_resp_bits_hx = ptw_resp_hx ; 
  assign  ptw_io_requestor_0_resp_bits_pte_ppn = ptw_r_pte_ppn ; 
  assign  ptw_io_requestor_0_resp_bits_pte_d = ptw_r_pte_d ; 
  assign  ptw_io_requestor_0_resp_bits_pte_a = ptw_r_pte_a ; 
  assign  ptw_io_requestor_0_resp_bits_pte_g = ptw_r_pte_g ; 
  assign  ptw_io_requestor_0_resp_bits_pte_u = ptw_r_pte_u ; 
  assign  ptw_io_requestor_0_resp_bits_pte_x = ptw_r_pte_x ; 
  assign  ptw_io_requestor_0_resp_bits_pte_w = ptw_r_pte_w ; 
  assign  ptw_io_requestor_0_resp_bits_pte_r = ptw_r_pte_r ; 
  assign  ptw_io_requestor_0_resp_bits_pte_v = ptw_r_pte_v ; 
  assign  ptw_io_requestor_0_resp_bits_gpa_is_pte =~ ptw_stage2_final ; 
  assign  ptw_io_requestor_0_status_debug = ptw_io_dpath_status_debug ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_l = ptw_io_dpath_pmp_0_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_a = ptw_io_dpath_pmp_0_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_x = ptw_io_dpath_pmp_0_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_w = ptw_io_dpath_pmp_0_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_r = ptw_io_dpath_pmp_0_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_0_addr = ptw_io_dpath_pmp_0_addr ; 
  assign  ptw_io_requestor_0_pmp_0_mask = ptw_io_dpath_pmp_0_mask ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_l = ptw_io_dpath_pmp_1_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_a = ptw_io_dpath_pmp_1_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_x = ptw_io_dpath_pmp_1_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_w = ptw_io_dpath_pmp_1_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_r = ptw_io_dpath_pmp_1_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_1_addr = ptw_io_dpath_pmp_1_addr ; 
  assign  ptw_io_requestor_0_pmp_1_mask = ptw_io_dpath_pmp_1_mask ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_l = ptw_io_dpath_pmp_2_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_a = ptw_io_dpath_pmp_2_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_x = ptw_io_dpath_pmp_2_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_w = ptw_io_dpath_pmp_2_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_r = ptw_io_dpath_pmp_2_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_2_addr = ptw_io_dpath_pmp_2_addr ; 
  assign  ptw_io_requestor_0_pmp_2_mask = ptw_io_dpath_pmp_2_mask ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_l = ptw_io_dpath_pmp_3_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_a = ptw_io_dpath_pmp_3_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_x = ptw_io_dpath_pmp_3_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_w = ptw_io_dpath_pmp_3_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_r = ptw_io_dpath_pmp_3_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_3_addr = ptw_io_dpath_pmp_3_addr ; 
  assign  ptw_io_requestor_0_pmp_3_mask = ptw_io_dpath_pmp_3_mask ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_l = ptw_io_dpath_pmp_4_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_a = ptw_io_dpath_pmp_4_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_x = ptw_io_dpath_pmp_4_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_w = ptw_io_dpath_pmp_4_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_r = ptw_io_dpath_pmp_4_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_4_addr = ptw_io_dpath_pmp_4_addr ; 
  assign  ptw_io_requestor_0_pmp_4_mask = ptw_io_dpath_pmp_4_mask ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_l = ptw_io_dpath_pmp_5_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_a = ptw_io_dpath_pmp_5_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_x = ptw_io_dpath_pmp_5_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_w = ptw_io_dpath_pmp_5_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_r = ptw_io_dpath_pmp_5_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_5_addr = ptw_io_dpath_pmp_5_addr ; 
  assign  ptw_io_requestor_0_pmp_5_mask = ptw_io_dpath_pmp_5_mask ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_l = ptw_io_dpath_pmp_6_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_a = ptw_io_dpath_pmp_6_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_x = ptw_io_dpath_pmp_6_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_w = ptw_io_dpath_pmp_6_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_r = ptw_io_dpath_pmp_6_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_6_addr = ptw_io_dpath_pmp_6_addr ; 
  assign  ptw_io_requestor_0_pmp_6_mask = ptw_io_dpath_pmp_6_mask ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_l = ptw_io_dpath_pmp_7_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_a = ptw_io_dpath_pmp_7_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_x = ptw_io_dpath_pmp_7_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_w = ptw_io_dpath_pmp_7_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_r = ptw_io_dpath_pmp_7_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_7_addr = ptw_io_dpath_pmp_7_addr ; 
  assign  ptw_io_requestor_0_pmp_7_mask = ptw_io_dpath_pmp_7_mask ; 
  assign  ptw_io_requestor_1_resp_bits_ae_ptw = ptw_resp_ae_ptw ; 
  assign  ptw_io_requestor_1_resp_bits_ae_final = ptw_resp_ae_final ; 
  assign  ptw_io_requestor_1_resp_bits_pf = ptw_resp_pf ; 
  assign  ptw_io_requestor_1_resp_bits_gf = ptw_resp_gf ; 
  assign  ptw_io_requestor_1_resp_bits_hr = ptw_resp_hr ; 
  assign  ptw_io_requestor_1_resp_bits_hw = ptw_resp_hw ; 
  assign  ptw_io_requestor_1_resp_bits_hx = ptw_resp_hx ; 
  assign  ptw_io_requestor_1_resp_bits_pte_ppn = ptw_r_pte_ppn ; 
  assign  ptw_io_requestor_1_resp_bits_pte_d = ptw_r_pte_d ; 
  assign  ptw_io_requestor_1_resp_bits_pte_a = ptw_r_pte_a ; 
  assign  ptw_io_requestor_1_resp_bits_pte_g = ptw_r_pte_g ; 
  assign  ptw_io_requestor_1_resp_bits_pte_u = ptw_r_pte_u ; 
  assign  ptw_io_requestor_1_resp_bits_pte_x = ptw_r_pte_x ; 
  assign  ptw_io_requestor_1_resp_bits_pte_w = ptw_r_pte_w ; 
  assign  ptw_io_requestor_1_resp_bits_pte_r = ptw_r_pte_r ; 
  assign  ptw_io_requestor_1_resp_bits_pte_v = ptw_r_pte_v ; 
  assign  ptw_io_requestor_1_resp_bits_gpa_is_pte =~ ptw_stage2_final ; 
  assign  ptw_io_requestor_1_status_debug = ptw_io_dpath_status_debug ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_l = ptw_io_dpath_pmp_0_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_a = ptw_io_dpath_pmp_0_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_x = ptw_io_dpath_pmp_0_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_w = ptw_io_dpath_pmp_0_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_r = ptw_io_dpath_pmp_0_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_0_addr = ptw_io_dpath_pmp_0_addr ; 
  assign  ptw_io_requestor_1_pmp_0_mask = ptw_io_dpath_pmp_0_mask ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_l = ptw_io_dpath_pmp_1_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_a = ptw_io_dpath_pmp_1_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_x = ptw_io_dpath_pmp_1_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_w = ptw_io_dpath_pmp_1_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_r = ptw_io_dpath_pmp_1_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_1_addr = ptw_io_dpath_pmp_1_addr ; 
  assign  ptw_io_requestor_1_pmp_1_mask = ptw_io_dpath_pmp_1_mask ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_l = ptw_io_dpath_pmp_2_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_a = ptw_io_dpath_pmp_2_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_x = ptw_io_dpath_pmp_2_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_w = ptw_io_dpath_pmp_2_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_r = ptw_io_dpath_pmp_2_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_2_addr = ptw_io_dpath_pmp_2_addr ; 
  assign  ptw_io_requestor_1_pmp_2_mask = ptw_io_dpath_pmp_2_mask ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_l = ptw_io_dpath_pmp_3_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_a = ptw_io_dpath_pmp_3_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_x = ptw_io_dpath_pmp_3_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_w = ptw_io_dpath_pmp_3_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_r = ptw_io_dpath_pmp_3_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_3_addr = ptw_io_dpath_pmp_3_addr ; 
  assign  ptw_io_requestor_1_pmp_3_mask = ptw_io_dpath_pmp_3_mask ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_l = ptw_io_dpath_pmp_4_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_a = ptw_io_dpath_pmp_4_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_x = ptw_io_dpath_pmp_4_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_w = ptw_io_dpath_pmp_4_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_r = ptw_io_dpath_pmp_4_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_4_addr = ptw_io_dpath_pmp_4_addr ; 
  assign  ptw_io_requestor_1_pmp_4_mask = ptw_io_dpath_pmp_4_mask ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_l = ptw_io_dpath_pmp_5_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_a = ptw_io_dpath_pmp_5_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_x = ptw_io_dpath_pmp_5_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_w = ptw_io_dpath_pmp_5_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_r = ptw_io_dpath_pmp_5_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_5_addr = ptw_io_dpath_pmp_5_addr ; 
  assign  ptw_io_requestor_1_pmp_5_mask = ptw_io_dpath_pmp_5_mask ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_l = ptw_io_dpath_pmp_6_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_a = ptw_io_dpath_pmp_6_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_x = ptw_io_dpath_pmp_6_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_w = ptw_io_dpath_pmp_6_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_r = ptw_io_dpath_pmp_6_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_6_addr = ptw_io_dpath_pmp_6_addr ; 
  assign  ptw_io_requestor_1_pmp_6_mask = ptw_io_dpath_pmp_6_mask ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_l = ptw_io_dpath_pmp_7_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_a = ptw_io_dpath_pmp_7_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_x = ptw_io_dpath_pmp_7_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_w = ptw_io_dpath_pmp_7_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_r = ptw_io_dpath_pmp_7_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_7_addr = ptw_io_dpath_pmp_7_addr ; 
  assign  ptw_io_requestor_1_pmp_7_mask = ptw_io_dpath_pmp_7_mask ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_0_value = ptw_io_dpath_customCSRs_csrs_0_value ;
    assign ptw_clock = clock;
    assign ptw_reset = reset;
    assign ptw_io_requestor_0_req_bits_bits_addr = _dcache_io_ptw_req_bits_bits_addr;
    assign ptw_io_requestor_0_req_bits_bits_need_gpa = _dcache_io_ptw_req_bits_bits_need_gpa;
    assign ptw_io_requestor_0_req_bits_bits_vstage1 = _dcache_io_ptw_req_bits_bits_vstage1;
    assign ptw_io_requestor_0_req_bits_bits_stage2 = _dcache_io_ptw_req_bits_bits_stage2;
    assign _ptw_io_requestor_0_resp_bits_ae_ptw = ptw_io_requestor_0_resp_bits_ae_ptw;
    assign _ptw_io_requestor_0_resp_bits_ae_final = ptw_io_requestor_0_resp_bits_ae_final;
    assign _ptw_io_requestor_0_resp_bits_pf = ptw_io_requestor_0_resp_bits_pf;
    assign _ptw_io_requestor_0_resp_bits_gf = ptw_io_requestor_0_resp_bits_gf;
    assign _ptw_io_requestor_0_resp_bits_hr = ptw_io_requestor_0_resp_bits_hr;
    assign _ptw_io_requestor_0_resp_bits_hw = ptw_io_requestor_0_resp_bits_hw;
    assign _ptw_io_requestor_0_resp_bits_hx = ptw_io_requestor_0_resp_bits_hx;
    assign _ptw_io_requestor_0_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn;
    assign _ptw_io_requestor_0_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d;
    assign _ptw_io_requestor_0_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a;
    assign _ptw_io_requestor_0_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g;
    assign _ptw_io_requestor_0_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u;
    assign _ptw_io_requestor_0_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x;
    assign _ptw_io_requestor_0_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w;
    assign _ptw_io_requestor_0_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r;
    assign _ptw_io_requestor_0_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v;
    assign _ptw_io_requestor_0_resp_bits_gpa_is_pte = ptw_io_requestor_0_resp_bits_gpa_is_pte;
    assign _ptw_io_requestor_0_status_debug = ptw_io_requestor_0_status_debug;
    assign _ptw_io_requestor_0_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l;
    assign _ptw_io_requestor_0_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a;
    assign _ptw_io_requestor_0_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x;
    assign _ptw_io_requestor_0_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w;
    assign _ptw_io_requestor_0_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r;
    assign _ptw_io_requestor_0_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr;
    assign _ptw_io_requestor_0_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask;
    assign _ptw_io_requestor_0_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l;
    assign _ptw_io_requestor_0_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a;
    assign _ptw_io_requestor_0_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x;
    assign _ptw_io_requestor_0_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w;
    assign _ptw_io_requestor_0_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r;
    assign _ptw_io_requestor_0_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr;
    assign _ptw_io_requestor_0_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask;
    assign _ptw_io_requestor_0_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l;
    assign _ptw_io_requestor_0_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a;
    assign _ptw_io_requestor_0_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x;
    assign _ptw_io_requestor_0_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w;
    assign _ptw_io_requestor_0_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r;
    assign _ptw_io_requestor_0_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr;
    assign _ptw_io_requestor_0_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask;
    assign _ptw_io_requestor_0_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l;
    assign _ptw_io_requestor_0_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a;
    assign _ptw_io_requestor_0_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x;
    assign _ptw_io_requestor_0_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w;
    assign _ptw_io_requestor_0_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r;
    assign _ptw_io_requestor_0_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr;
    assign _ptw_io_requestor_0_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask;
    assign _ptw_io_requestor_0_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l;
    assign _ptw_io_requestor_0_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a;
    assign _ptw_io_requestor_0_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x;
    assign _ptw_io_requestor_0_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w;
    assign _ptw_io_requestor_0_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r;
    assign _ptw_io_requestor_0_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr;
    assign _ptw_io_requestor_0_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask;
    assign _ptw_io_requestor_0_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l;
    assign _ptw_io_requestor_0_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a;
    assign _ptw_io_requestor_0_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x;
    assign _ptw_io_requestor_0_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w;
    assign _ptw_io_requestor_0_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r;
    assign _ptw_io_requestor_0_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr;
    assign _ptw_io_requestor_0_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask;
    assign _ptw_io_requestor_0_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l;
    assign _ptw_io_requestor_0_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a;
    assign _ptw_io_requestor_0_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x;
    assign _ptw_io_requestor_0_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w;
    assign _ptw_io_requestor_0_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r;
    assign _ptw_io_requestor_0_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr;
    assign _ptw_io_requestor_0_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask;
    assign _ptw_io_requestor_0_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l;
    assign _ptw_io_requestor_0_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a;
    assign _ptw_io_requestor_0_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x;
    assign _ptw_io_requestor_0_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w;
    assign _ptw_io_requestor_0_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r;
    assign _ptw_io_requestor_0_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr;
    assign _ptw_io_requestor_0_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask;
    assign ptw_io_requestor_1_req_bits_valid = _frontend_io_ptw_req_bits_valid;
    assign ptw_io_requestor_1_req_bits_bits_addr = _frontend_io_ptw_req_bits_bits_addr;
    assign ptw_io_requestor_1_req_bits_bits_need_gpa = _frontend_io_ptw_req_bits_bits_need_gpa;
    assign ptw_io_requestor_1_req_bits_bits_vstage1 = _frontend_io_ptw_req_bits_bits_vstage1;
    assign ptw_io_requestor_1_req_bits_bits_stage2 = _frontend_io_ptw_req_bits_bits_stage2;
    assign _ptw_io_requestor_1_resp_bits_ae_ptw = ptw_io_requestor_1_resp_bits_ae_ptw;
    assign _ptw_io_requestor_1_resp_bits_ae_final = ptw_io_requestor_1_resp_bits_ae_final;
    assign _ptw_io_requestor_1_resp_bits_pf = ptw_io_requestor_1_resp_bits_pf;
    assign _ptw_io_requestor_1_resp_bits_gf = ptw_io_requestor_1_resp_bits_gf;
    assign _ptw_io_requestor_1_resp_bits_hr = ptw_io_requestor_1_resp_bits_hr;
    assign _ptw_io_requestor_1_resp_bits_hw = ptw_io_requestor_1_resp_bits_hw;
    assign _ptw_io_requestor_1_resp_bits_hx = ptw_io_requestor_1_resp_bits_hx;
    assign _ptw_io_requestor_1_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn;
    assign _ptw_io_requestor_1_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d;
    assign _ptw_io_requestor_1_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a;
    assign _ptw_io_requestor_1_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g;
    assign _ptw_io_requestor_1_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u;
    assign _ptw_io_requestor_1_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x;
    assign _ptw_io_requestor_1_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w;
    assign _ptw_io_requestor_1_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r;
    assign _ptw_io_requestor_1_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v;
    assign _ptw_io_requestor_1_resp_bits_gpa_is_pte = ptw_io_requestor_1_resp_bits_gpa_is_pte;
    assign _ptw_io_requestor_1_status_debug = ptw_io_requestor_1_status_debug;
    assign _ptw_io_requestor_1_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l;
    assign _ptw_io_requestor_1_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a;
    assign _ptw_io_requestor_1_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x;
    assign _ptw_io_requestor_1_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w;
    assign _ptw_io_requestor_1_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r;
    assign _ptw_io_requestor_1_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr;
    assign _ptw_io_requestor_1_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask;
    assign _ptw_io_requestor_1_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l;
    assign _ptw_io_requestor_1_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a;
    assign _ptw_io_requestor_1_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x;
    assign _ptw_io_requestor_1_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w;
    assign _ptw_io_requestor_1_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r;
    assign _ptw_io_requestor_1_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr;
    assign _ptw_io_requestor_1_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask;
    assign _ptw_io_requestor_1_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l;
    assign _ptw_io_requestor_1_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a;
    assign _ptw_io_requestor_1_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x;
    assign _ptw_io_requestor_1_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w;
    assign _ptw_io_requestor_1_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r;
    assign _ptw_io_requestor_1_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr;
    assign _ptw_io_requestor_1_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask;
    assign _ptw_io_requestor_1_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l;
    assign _ptw_io_requestor_1_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a;
    assign _ptw_io_requestor_1_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x;
    assign _ptw_io_requestor_1_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w;
    assign _ptw_io_requestor_1_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r;
    assign _ptw_io_requestor_1_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr;
    assign _ptw_io_requestor_1_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask;
    assign _ptw_io_requestor_1_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l;
    assign _ptw_io_requestor_1_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a;
    assign _ptw_io_requestor_1_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x;
    assign _ptw_io_requestor_1_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w;
    assign _ptw_io_requestor_1_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r;
    assign _ptw_io_requestor_1_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr;
    assign _ptw_io_requestor_1_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask;
    assign _ptw_io_requestor_1_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l;
    assign _ptw_io_requestor_1_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a;
    assign _ptw_io_requestor_1_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x;
    assign _ptw_io_requestor_1_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w;
    assign _ptw_io_requestor_1_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r;
    assign _ptw_io_requestor_1_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr;
    assign _ptw_io_requestor_1_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask;
    assign _ptw_io_requestor_1_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l;
    assign _ptw_io_requestor_1_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a;
    assign _ptw_io_requestor_1_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x;
    assign _ptw_io_requestor_1_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w;
    assign _ptw_io_requestor_1_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r;
    assign _ptw_io_requestor_1_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr;
    assign _ptw_io_requestor_1_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask;
    assign _ptw_io_requestor_1_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l;
    assign _ptw_io_requestor_1_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a;
    assign _ptw_io_requestor_1_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x;
    assign _ptw_io_requestor_1_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w;
    assign _ptw_io_requestor_1_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r;
    assign _ptw_io_requestor_1_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr;
    assign _ptw_io_requestor_1_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask;
    assign _ptw_io_requestor_1_customCSRs_csrs_0_value = ptw_io_requestor_1_customCSRs_csrs_0_value;
    assign ptw_io_dpath_sfence_valid = _core_io_ptw_sfence_valid;
    assign ptw_io_dpath_sfence_bits_rs1 = _core_io_ptw_sfence_bits_rs1;
    assign ptw_io_dpath_status_debug = _core_io_ptw_status_debug;
    assign ptw_io_dpath_pmp_0_cfg_l = _core_io_ptw_pmp_0_cfg_l;
    assign ptw_io_dpath_pmp_0_cfg_a = _core_io_ptw_pmp_0_cfg_a;
    assign ptw_io_dpath_pmp_0_cfg_x = _core_io_ptw_pmp_0_cfg_x;
    assign ptw_io_dpath_pmp_0_cfg_w = _core_io_ptw_pmp_0_cfg_w;
    assign ptw_io_dpath_pmp_0_cfg_r = _core_io_ptw_pmp_0_cfg_r;
    assign ptw_io_dpath_pmp_0_addr = _core_io_ptw_pmp_0_addr;
    assign ptw_io_dpath_pmp_0_mask = _core_io_ptw_pmp_0_mask;
    assign ptw_io_dpath_pmp_1_cfg_l = _core_io_ptw_pmp_1_cfg_l;
    assign ptw_io_dpath_pmp_1_cfg_a = _core_io_ptw_pmp_1_cfg_a;
    assign ptw_io_dpath_pmp_1_cfg_x = _core_io_ptw_pmp_1_cfg_x;
    assign ptw_io_dpath_pmp_1_cfg_w = _core_io_ptw_pmp_1_cfg_w;
    assign ptw_io_dpath_pmp_1_cfg_r = _core_io_ptw_pmp_1_cfg_r;
    assign ptw_io_dpath_pmp_1_addr = _core_io_ptw_pmp_1_addr;
    assign ptw_io_dpath_pmp_1_mask = _core_io_ptw_pmp_1_mask;
    assign ptw_io_dpath_pmp_2_cfg_l = _core_io_ptw_pmp_2_cfg_l;
    assign ptw_io_dpath_pmp_2_cfg_a = _core_io_ptw_pmp_2_cfg_a;
    assign ptw_io_dpath_pmp_2_cfg_x = _core_io_ptw_pmp_2_cfg_x;
    assign ptw_io_dpath_pmp_2_cfg_w = _core_io_ptw_pmp_2_cfg_w;
    assign ptw_io_dpath_pmp_2_cfg_r = _core_io_ptw_pmp_2_cfg_r;
    assign ptw_io_dpath_pmp_2_addr = _core_io_ptw_pmp_2_addr;
    assign ptw_io_dpath_pmp_2_mask = _core_io_ptw_pmp_2_mask;
    assign ptw_io_dpath_pmp_3_cfg_l = _core_io_ptw_pmp_3_cfg_l;
    assign ptw_io_dpath_pmp_3_cfg_a = _core_io_ptw_pmp_3_cfg_a;
    assign ptw_io_dpath_pmp_3_cfg_x = _core_io_ptw_pmp_3_cfg_x;
    assign ptw_io_dpath_pmp_3_cfg_w = _core_io_ptw_pmp_3_cfg_w;
    assign ptw_io_dpath_pmp_3_cfg_r = _core_io_ptw_pmp_3_cfg_r;
    assign ptw_io_dpath_pmp_3_addr = _core_io_ptw_pmp_3_addr;
    assign ptw_io_dpath_pmp_3_mask = _core_io_ptw_pmp_3_mask;
    assign ptw_io_dpath_pmp_4_cfg_l = _core_io_ptw_pmp_4_cfg_l;
    assign ptw_io_dpath_pmp_4_cfg_a = _core_io_ptw_pmp_4_cfg_a;
    assign ptw_io_dpath_pmp_4_cfg_x = _core_io_ptw_pmp_4_cfg_x;
    assign ptw_io_dpath_pmp_4_cfg_w = _core_io_ptw_pmp_4_cfg_w;
    assign ptw_io_dpath_pmp_4_cfg_r = _core_io_ptw_pmp_4_cfg_r;
    assign ptw_io_dpath_pmp_4_addr = _core_io_ptw_pmp_4_addr;
    assign ptw_io_dpath_pmp_4_mask = _core_io_ptw_pmp_4_mask;
    assign ptw_io_dpath_pmp_5_cfg_l = _core_io_ptw_pmp_5_cfg_l;
    assign ptw_io_dpath_pmp_5_cfg_a = _core_io_ptw_pmp_5_cfg_a;
    assign ptw_io_dpath_pmp_5_cfg_x = _core_io_ptw_pmp_5_cfg_x;
    assign ptw_io_dpath_pmp_5_cfg_w = _core_io_ptw_pmp_5_cfg_w;
    assign ptw_io_dpath_pmp_5_cfg_r = _core_io_ptw_pmp_5_cfg_r;
    assign ptw_io_dpath_pmp_5_addr = _core_io_ptw_pmp_5_addr;
    assign ptw_io_dpath_pmp_5_mask = _core_io_ptw_pmp_5_mask;
    assign ptw_io_dpath_pmp_6_cfg_l = _core_io_ptw_pmp_6_cfg_l;
    assign ptw_io_dpath_pmp_6_cfg_a = _core_io_ptw_pmp_6_cfg_a;
    assign ptw_io_dpath_pmp_6_cfg_x = _core_io_ptw_pmp_6_cfg_x;
    assign ptw_io_dpath_pmp_6_cfg_w = _core_io_ptw_pmp_6_cfg_w;
    assign ptw_io_dpath_pmp_6_cfg_r = _core_io_ptw_pmp_6_cfg_r;
    assign ptw_io_dpath_pmp_6_addr = _core_io_ptw_pmp_6_addr;
    assign ptw_io_dpath_pmp_6_mask = _core_io_ptw_pmp_6_mask;
    assign ptw_io_dpath_pmp_7_cfg_l = _core_io_ptw_pmp_7_cfg_l;
    assign ptw_io_dpath_pmp_7_cfg_a = _core_io_ptw_pmp_7_cfg_a;
    assign ptw_io_dpath_pmp_7_cfg_x = _core_io_ptw_pmp_7_cfg_x;
    assign ptw_io_dpath_pmp_7_cfg_w = _core_io_ptw_pmp_7_cfg_w;
    assign ptw_io_dpath_pmp_7_cfg_r = _core_io_ptw_pmp_7_cfg_r;
    assign ptw_io_dpath_pmp_7_addr = _core_io_ptw_pmp_7_addr;
    assign ptw_io_dpath_pmp_7_mask = _core_io_ptw_pmp_7_mask;
    assign ptw_io_dpath_customCSRs_csrs_0_value = _core_io_ptw_customCSRs_csrs_0_value;
    
  wire core_clock;
    wire core_reset;
    wire core_io_hartid;
    wire core_io_interrupts_debug;
    wire core_io_interrupts_mtip;
    wire core_io_interrupts_msip;
    wire core_io_interrupts_meip;
    wire core_io_imem_might_request;
    wire core_io_imem_req_valid;
    wire[31:0] core_io_imem_req_bits_pc;
    wire core_io_imem_req_bits_speculative;
    wire core_io_imem_sfence_valid;
    wire core_io_imem_resp_ready;
    wire core_io_imem_resp_valid;
    wire[1:0] core_io_imem_resp_bits_btb_cfiType;
    wire core_io_imem_resp_bits_btb_taken;
    wire[1:0] core_io_imem_resp_bits_btb_mask;
    wire core_io_imem_resp_bits_btb_bridx;
    wire[31:0] core_io_imem_resp_bits_btb_target;
    wire core_io_imem_resp_bits_btb_entry;
    wire[7:0] core_io_imem_resp_bits_btb_bht_history;
    wire core_io_imem_resp_bits_btb_bht_value;
    wire[31:0] core_io_imem_resp_bits_pc;
    wire[31:0] core_io_imem_resp_bits_data;
    wire[1:0] core_io_imem_resp_bits_mask;
    wire core_io_imem_resp_bits_xcpt_pf_inst;
    wire core_io_imem_resp_bits_xcpt_gf_inst;
    wire core_io_imem_resp_bits_xcpt_ae_inst;
    wire core_io_imem_resp_bits_replay;
    wire core_io_imem_gpa_valid;
    wire[31:0] core_io_imem_gpa_bits;
    wire core_io_imem_btb_update_valid;
    wire core_io_imem_bht_update_valid;
    wire core_io_imem_flush_icache;
    wire core_io_imem_progress;
    wire core_io_dmem_req_ready;
    wire core_io_dmem_req_valid;
    wire[31:0] core_io_dmem_req_bits_addr;
    wire[6:0] core_io_dmem_req_bits_tag;
    wire[4:0] core_io_dmem_req_bits_cmd;
    wire[1:0] core_io_dmem_req_bits_size;
    wire core_io_dmem_req_bits_signed;
    wire core_io_dmem_req_bits_dv;
    wire core_io_dmem_s1_kill;
    wire[31:0] core_io_dmem_s1_data_data;
    wire core_io_dmem_s2_nack;
    wire core_io_dmem_resp_valid;
    wire[6:0] core_io_dmem_resp_bits_tag;
    wire[31:0] core_io_dmem_resp_bits_data;
    wire core_io_dmem_resp_bits_replay;
    wire core_io_dmem_resp_bits_has_data;
    wire[31:0] core_io_dmem_resp_bits_data_word_bypass;
    wire core_io_dmem_replay_next;
    wire core_io_dmem_s2_xcpt_ma_ld;
    wire core_io_dmem_s2_xcpt_ma_st;
    wire core_io_dmem_s2_xcpt_pf_ld;
    wire core_io_dmem_s2_xcpt_pf_st;
    wire core_io_dmem_s2_xcpt_ae_ld;
    wire core_io_dmem_s2_xcpt_ae_st;
    wire core_io_dmem_ordered;
    wire core_io_dmem_perf_grant;
    wire core_io_ptw_sfence_valid;
    wire core_io_ptw_sfence_bits_rs1;
    wire core_io_ptw_status_debug;
    wire core_io_ptw_pmp_0_cfg_l;
    wire[1:0] core_io_ptw_pmp_0_cfg_a;
    wire core_io_ptw_pmp_0_cfg_x;
    wire core_io_ptw_pmp_0_cfg_w;
    wire core_io_ptw_pmp_0_cfg_r;
    wire[29:0] core_io_ptw_pmp_0_addr;
    wire[31:0] core_io_ptw_pmp_0_mask;
    wire core_io_ptw_pmp_1_cfg_l;
    wire[1:0] core_io_ptw_pmp_1_cfg_a;
    wire core_io_ptw_pmp_1_cfg_x;
    wire core_io_ptw_pmp_1_cfg_w;
    wire core_io_ptw_pmp_1_cfg_r;
    wire[29:0] core_io_ptw_pmp_1_addr;
    wire[31:0] core_io_ptw_pmp_1_mask;
    wire core_io_ptw_pmp_2_cfg_l;
    wire[1:0] core_io_ptw_pmp_2_cfg_a;
    wire core_io_ptw_pmp_2_cfg_x;
    wire core_io_ptw_pmp_2_cfg_w;
    wire core_io_ptw_pmp_2_cfg_r;
    wire[29:0] core_io_ptw_pmp_2_addr;
    wire[31:0] core_io_ptw_pmp_2_mask;
    wire core_io_ptw_pmp_3_cfg_l;
    wire[1:0] core_io_ptw_pmp_3_cfg_a;
    wire core_io_ptw_pmp_3_cfg_x;
    wire core_io_ptw_pmp_3_cfg_w;
    wire core_io_ptw_pmp_3_cfg_r;
    wire[29:0] core_io_ptw_pmp_3_addr;
    wire[31:0] core_io_ptw_pmp_3_mask;
    wire core_io_ptw_pmp_4_cfg_l;
    wire[1:0] core_io_ptw_pmp_4_cfg_a;
    wire core_io_ptw_pmp_4_cfg_x;
    wire core_io_ptw_pmp_4_cfg_w;
    wire core_io_ptw_pmp_4_cfg_r;
    wire[29:0] core_io_ptw_pmp_4_addr;
    wire[31:0] core_io_ptw_pmp_4_mask;
    wire core_io_ptw_pmp_5_cfg_l;
    wire[1:0] core_io_ptw_pmp_5_cfg_a;
    wire core_io_ptw_pmp_5_cfg_x;
    wire core_io_ptw_pmp_5_cfg_w;
    wire core_io_ptw_pmp_5_cfg_r;
    wire[29:0] core_io_ptw_pmp_5_addr;
    wire[31:0] core_io_ptw_pmp_5_mask;
    wire core_io_ptw_pmp_6_cfg_l;
    wire[1:0] core_io_ptw_pmp_6_cfg_a;
    wire core_io_ptw_pmp_6_cfg_x;
    wire core_io_ptw_pmp_6_cfg_w;
    wire core_io_ptw_pmp_6_cfg_r;
    wire[29:0] core_io_ptw_pmp_6_addr;
    wire[31:0] core_io_ptw_pmp_6_mask;
    wire core_io_ptw_pmp_7_cfg_l;
    wire[1:0] core_io_ptw_pmp_7_cfg_a;
    wire core_io_ptw_pmp_7_cfg_x;
    wire core_io_ptw_pmp_7_cfg_w;
    wire core_io_ptw_pmp_7_cfg_r;
    wire[29:0] core_io_ptw_pmp_7_addr;
    wire[31:0] core_io_ptw_pmp_7_mask;
    wire[31:0] core_io_ptw_customCSRs_csrs_0_value;
    wire core_io_trace_insns_0_valid;
    wire[31:0] core_io_trace_insns_0_iaddr;
    wire[31:0] core_io_trace_insns_0_insn;
    wire[2:0] core_io_trace_insns_0_priv;
    wire core_io_trace_insns_0_exception;
    wire core_io_trace_insns_0_interrupt;
    wire[31:0] core_io_trace_insns_0_cause;
    wire[31:0] core_io_trace_insns_0_tval;
    wire[63:0] core_io_trace_time;
    wire core_io_bpwatch_0_valid_0;
    wire[2:0] core_io_bpwatch_0_action;
    wire core_io_wfi;

    wire[4:0] core_id_raddr3 ; 
    wire core__io_dmem_req_valid_output ; 
    wire core__GEN ; 
    wire core__div_io_req_ready ; 
    wire core__div_io_resp_valid ; 
    wire[4:0] core__div_io_resp_bits_tag ; 
    wire[31:0] core__alu_io_out ; 
    wire core__alu_io_cmp_out ; 
    wire core__bpu_io_xcpt_if ; 
    wire core__bpu_io_xcpt_ld ; 
    wire core__bpu_io_xcpt_st ; 
    wire core__bpu_io_debug_if ; 
    wire core__bpu_io_debug_ld ; 
    wire core__bpu_io_debug_st ; 
    wire core__bpu_io_bpwatch_0_rvalid_0 ; 
    wire core__bpu_io_bpwatch_0_wvalid_0 ; 
    wire core__bpu_io_bpwatch_0_ivalid_0 ; 
    wire[31:0] core__csr_io_rw_rdata ; 
    wire core__csr_io_decode_0_read_illegal ; 
    wire core__csr_io_decode_0_write_illegal ; 
    wire core__csr_io_decode_0_write_flush ; 
    wire core__csr_io_decode_0_system_illegal ; 
    wire core__csr_io_decode_0_virtual_access_illegal ; 
    wire core__csr_io_decode_0_virtual_system_illegal ; 
    wire core__csr_io_csr_stall ; 
    wire core__csr_io_eret ; 
    wire core__csr_io_singleStep ; 
    wire core__csr_io_status_debug ; 
    wire[31:0] core__csr_io_status_isa ; 
    wire core__csr_io_status_dv ; 
    wire core__csr_io_status_v ; 
    wire[31:0] core__csr_io_evec ; 
    wire[31:0] core__csr_io_time ; 
    wire core__csr_io_interrupt ; 
    wire[31:0] core__csr_io_interrupt_cause ; 
    wire core__csr_io_bp_0_control_action ; 
    wire[1:0] core__csr_io_bp_0_control_tmatch ; 
    wire core__csr_io_bp_0_control_x ; 
    wire core__csr_io_bp_0_control_w ; 
    wire core__csr_io_bp_0_control_r ; 
    wire[31:0] core__csr_io_bp_0_address ; 
    wire core__csr_io_inhibit_cycle ; 
    wire core__csr_io_trace_0_valid ; 
    wire[31:0] core__csr_io_trace_0_iaddr ; 
    wire[31:0] core__csr_io_trace_0_insn ; 
    wire[2:0] core__csr_io_trace_0_priv ; 
    wire core__csr_io_trace_0_exception ; 
    wire[31:0] core__csr_io_customCSRs_0_value ; 
    wire[31:0] core__rf_ext_R0_data ; 
    wire[31:0] core__rf_ext_R1_data ; 
    wire[31:0] core__ibuf_io_pc ; 
    wire[1:0] core__ibuf_io_btb_resp_cfiType ; 
    wire core__ibuf_io_btb_resp_taken ; 
    wire[1:0] core__ibuf_io_btb_resp_mask ; 
    wire core__ibuf_io_btb_resp_bridx ; 
    wire[31:0] core__ibuf_io_btb_resp_target ; 
    wire core__ibuf_io_btb_resp_entry ; 
    wire[7:0] core__ibuf_io_btb_resp_bht_history ; 
    wire core__ibuf_io_btb_resp_bht_value ; 
    wire core__ibuf_io_inst_0_valid ; 
    wire core__ibuf_io_inst_0_bits_xcpt0_pf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt0_gf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt0_ae_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt1_pf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt1_gf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt1_ae_inst ; 
    wire core__ibuf_io_inst_0_bits_replay ; 
    wire core__ibuf_io_inst_0_bits_rvc ; 
    wire[31:0] core__ibuf_io_inst_0_bits_inst_bits ; 
    wire[4:0] core__ibuf_io_inst_0_bits_inst_rs1 ; 
    wire[31:0] core__ibuf_io_inst_0_bits_raw ; 
    wire[31:0] core_dcache_bypass_data = core_io_dmem_resp_bits_data_word_bypass ; 
    wire core_coreMonitorBundle_clock = core_clock ; 
    wire core_coreMonitorBundle_reset = core_reset ; 
    wire core_xrfWriteBundle_clock = core_clock ; 
    wire core_xrfWriteBundle_reset = core_reset ; 
    wire core_clock_en =1'h1; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_lo =2'h0; 
    wire core_hits_0 =1'h0; 
    wire core_hits_1 =1'h0; 
    wire core_hits_2 =1'h0; 
    wire core_hits_3 =1'h0; 
    wire core_hits_4 =1'h0; 
    wire core_hits_5 =1'h0; 
    wire core_hits_6 =1'h0; 
    wire core_hits_7 =1'h0; 
    wire core_hits_8 =1'h0; 
    wire core_hits_9 =1'h0; 
    wire core_hits_10 =1'h0; 
    wire core_hits_1_0 =1'h0; 
    wire core_hits_1_1 =1'h0; 
    wire core_hits_1_2 =1'h0; 
    wire core_hits_1_3 =1'h0; 
    wire core_hits_1_4 =1'h0; 
    wire core_hits_1_5 =1'h0; 
    wire core_hits_1_6 =1'h0; 
    wire core_hits_1_7 =1'h0; 
    wire core_hits_1_8 =1'h0; 
    wire core_hits_1_9 =1'h0; 
    wire core_hits_2_0 =1'h0; 
    wire core_hits_2_1 =1'h0; 
    wire core_hits_2_2 =1'h0; 
    wire core_hits_2_3 =1'h0; 
    wire core_hits_2_4 =1'h0; 
    wire core_hits_2_5 =1'h0; 
    wire core_id_npc_b0 =1'h0; 
    wire core_id_rocc_busy =1'h0; 
    wire core_ex_sfence =1'h0; 
    wire core_mem_br_target_b0 =1'h0; 
    wire core_mem_br_target_b0_1 =1'h0; 
    wire core_fpu_kill_mem =1'h0; 
    wire core_replay_wb_csr =1'h0; 
    wire core_csr_io_htval_htval_valid_dmem =1'h0; 
    wire core_fp_data_hazard_ex =1'h0; 
    wire core_fp_data_hazard_mem =1'h0; 
    wire core_fp_data_hazard_wb =1'h0; 
    wire core_coreMonitorBundle_wrenf =1'h0; 
    wire core_xrfWriteBundle_excpt =1'h0; 
    wire core_xrfWriteBundle_valid =1'h0; 
    wire core_xrfWriteBundle_wrenf =1'h0; 
    wire[31:0] core_csr_io_htval_htval_dmem =32'h0; 
    wire[31:0] core_xrfWriteBundle_pc =32'h0; 
    wire[31:0] core_xrfWriteBundle_rd0val =32'h0; 
    wire[31:0] core_xrfWriteBundle_rd1val =32'h0; 
    wire[31:0] core_xrfWriteBundle_inst =32'h0; 
    wire[4:0] core_xrfWriteBundle_rd0src =5'h0; 
    wire[4:0] core_xrfWriteBundle_rd1src =5'h0; 
    reg core_id_reg_pause ; 
    reg core_imem_might_request_reg ; 
    reg core_ex_ctrl_legal ; 
    reg core_ex_ctrl_fp ; 
    reg core_ex_ctrl_rocc ; 
    reg core_ex_ctrl_branch ; 
    reg core_ex_ctrl_jal ; 
    reg core_ex_ctrl_jalr ; 
    reg core_ex_ctrl_rxs2 ; 
    reg core_ex_ctrl_rxs1 ; reg[1:0] core_ex_ctrl_sel_alu2 ; reg[1:0] core_ex_ctrl_sel_alu1 ; reg[2:0] core_ex_ctrl_sel_imm ; 
    reg core_ex_ctrl_alu_dw ; reg[3:0] core_ex_ctrl_alu_fn ; 
    reg core_ex_ctrl_mem ; reg[4:0] core_ex_ctrl_mem_cmd ; 
    reg core_ex_ctrl_rfs1 ; 
    reg core_ex_ctrl_rfs2 ; 
    reg core_ex_ctrl_rfs3 ; 
    reg core_ex_ctrl_wfd ; 
    reg core_ex_ctrl_mul ; 
    reg core_ex_ctrl_div ; 
    reg core_ex_ctrl_wxd ; reg[2:0] core_ex_ctrl_csr ; 
    reg core_ex_ctrl_fence_i ; 
    reg core_ex_ctrl_fence ; 
    reg core_ex_ctrl_amo ; 
    reg core_ex_ctrl_dp ; 
    reg core_mem_ctrl_legal ; 
    reg core_mem_ctrl_fp ; 
    reg core_mem_ctrl_rocc ; 
    reg core_mem_ctrl_branch ; 
    reg core_mem_ctrl_jal ; 
    reg core_mem_ctrl_jalr ; 
    reg core_mem_ctrl_rxs2 ; 
    reg core_mem_ctrl_rxs1 ; reg[1:0] core_mem_ctrl_sel_alu2 ; reg[1:0] core_mem_ctrl_sel_alu1 ; reg[2:0] core_mem_ctrl_sel_imm ; 
    reg core_mem_ctrl_alu_dw ; reg[3:0] core_mem_ctrl_alu_fn ; 
    reg core_mem_ctrl_mem ; reg[4:0] core_mem_ctrl_mem_cmd ; 
    reg core_mem_ctrl_rfs1 ; 
    reg core_mem_ctrl_rfs2 ; 
    reg core_mem_ctrl_rfs3 ; 
    reg core_mem_ctrl_wfd ; 
    reg core_mem_ctrl_mul ; 
    reg core_mem_ctrl_div ; 
    reg core_mem_ctrl_wxd ; reg[2:0] core_mem_ctrl_csr ; 
    reg core_mem_ctrl_fence_i ; 
    reg core_mem_ctrl_fence ; 
    reg core_mem_ctrl_amo ; 
    reg core_mem_ctrl_dp ; 
    reg core_wb_ctrl_legal ; 
    reg core_wb_ctrl_fp ; 
    reg core_wb_ctrl_rocc ; 
    reg core_wb_ctrl_branch ; 
    reg core_wb_ctrl_jal ; 
    reg core_wb_ctrl_jalr ; 
    reg core_wb_ctrl_rxs2 ; 
    reg core_wb_ctrl_rxs1 ; reg[1:0] core_wb_ctrl_sel_alu2 ; reg[1:0] core_wb_ctrl_sel_alu1 ; reg[2:0] core_wb_ctrl_sel_imm ; 
    reg core_wb_ctrl_alu_dw ; reg[3:0] core_wb_ctrl_alu_fn ; 
    reg core_wb_ctrl_mem ; reg[4:0] core_wb_ctrl_mem_cmd ; 
    reg core_wb_ctrl_rfs1 ; 
    reg core_wb_ctrl_rfs2 ; 
    reg core_wb_ctrl_rfs3 ; 
    reg core_wb_ctrl_wfd ; 
    reg core_wb_ctrl_mul ; 
    reg core_wb_ctrl_div ; 
    reg core_wb_ctrl_wxd ; reg[2:0] core_wb_ctrl_csr ; 
    reg core_wb_ctrl_fence_i ; 
    reg core_wb_ctrl_fence ; 
    reg core_wb_ctrl_amo ; 
    reg core_wb_ctrl_dp ; 
    reg core_ex_reg_xcpt_interrupt ; 
    reg core_ex_reg_valid ; 
    reg core_ex_reg_rvc ; reg[1:0] core_ex_reg_btb_resp_cfiType ; 
    reg core_ex_reg_btb_resp_taken ; reg[1:0] core_ex_reg_btb_resp_mask ; 
    reg core_ex_reg_btb_resp_bridx ; reg[31:0] core_ex_reg_btb_resp_target ; 
    reg core_ex_reg_btb_resp_entry ; reg[7:0] core_ex_reg_btb_resp_bht_history ; 
    reg core_ex_reg_btb_resp_bht_value ; 
    reg core_ex_reg_xcpt ; 
    reg core_ex_reg_flush_pipe ; 
    reg core_ex_reg_load_use ; reg[31:0] core_ex_reg_cause ; 
    reg core_ex_reg_replay ; reg[31:0] core_ex_reg_pc ; reg[1:0] core_ex_reg_mem_size ; reg[31:0] core_ex_reg_inst ; reg[31:0] core_ex_reg_raw_inst ; 
    reg core_ex_reg_wphit_0 ; 
    reg core_mem_reg_xcpt_interrupt ; 
    reg core_mem_reg_valid ; 
    reg core_mem_reg_rvc ; reg[1:0] core_mem_reg_btb_resp_cfiType ; 
    reg core_mem_reg_btb_resp_taken ; reg[1:0] core_mem_reg_btb_resp_mask ; 
    reg core_mem_reg_btb_resp_bridx ; reg[31:0] core_mem_reg_btb_resp_target ; 
    reg core_mem_reg_btb_resp_entry ; reg[7:0] core_mem_reg_btb_resp_bht_history ; 
    reg core_mem_reg_btb_resp_bht_value ; 
    reg core_mem_reg_xcpt ; 
    reg core_mem_reg_replay ; 
    reg core_mem_reg_flush_pipe ; reg[31:0] core_mem_reg_cause ; 
    reg core_mem_reg_slow_bypass ; 
    wire core_mem_mem_cmd_bh = core_mem_reg_slow_bypass ; 
    reg core_mem_reg_load ; 
    reg core_mem_reg_store ; reg[31:0] core_mem_reg_pc ; reg[31:0] core_mem_reg_inst ; reg[1:0] core_mem_reg_mem_size ; 
    reg core_mem_reg_hls_or_dv ; reg[31:0] core_mem_reg_raw_inst ; reg[31:0] core_mem_reg_wdata ; reg[31:0] core_mem_reg_rs2 ; 
    reg core_mem_br_taken ; 
    reg core_mem_reg_wphit_0 ; 
    reg core_wb_reg_valid ; 
    reg core_wb_reg_xcpt ; 
    reg core_wb_reg_replay ; 
    reg core_wb_reg_flush_pipe ; reg[31:0] core_wb_reg_cause ; 
    reg core_wb_reg_sfence ; reg[31:0] core_wb_reg_pc ; reg[1:0] core_wb_reg_mem_size ; 
    reg core_wb_reg_hls_or_dv ; 
    reg core_wb_reg_hfence_v ; 
    reg core_wb_reg_hfence_g ; reg[31:0] core_wb_reg_inst ; reg[31:0] core_wb_reg_raw_inst ; reg[31:0] core_wb_reg_wdata ; reg[31:0] core_wb_reg_rs2 ; 
    reg core_wb_reg_wphit_0 ; 
    wire core_take_pc_mem ; 
    wire core_take_pc_wb ; 
    wire core_take_pc_mem_wb = core_take_pc_wb | core_take_pc_mem ; 
    wire core_id_ctrl_decoder_0 ; 
    wire core_id_ctrl_decoder_1 ; 
    wire core_id_ctrl_decoder_2 ; 
    wire core_id_ctrl_decoder_3 ; 
    wire core_id_ctrl_decoder_4 ; 
    wire core_id_ctrl_decoder_5 ; 
    wire core_id_ctrl_decoder_6 ; 
    wire core_id_ctrl_decoder_7 ; 
    wire[1:0] core_id_ctrl_decoder_8 ; 
    wire[1:0] core_id_ctrl_decoder_9 ; 
    wire[2:0] core_id_ctrl_decoder_10 ; 
    wire core_id_ctrl_decoder_11 ; 
    wire[3:0] core_id_ctrl_decoder_12 ; 
    wire core_id_ctrl_decoder_13 ; 
    wire[4:0] core_id_ctrl_decoder_14 ; 
    wire core_id_ctrl_decoder_15 ; 
    wire core_id_ctrl_decoder_16 ; 
    wire core_id_ctrl_decoder_17 ; 
    wire core_id_ctrl_decoder_18 ; 
    wire core_id_ctrl_decoder_19 ; 
    wire core_id_ctrl_decoder_20 ; 
    wire core_id_ctrl_decoder_21 ; 
    wire[2:0] core_id_ctrl_decoder_22 ; 
    wire core_id_ctrl_decoder_23 ; 
    wire core_id_ctrl_decoder_24 ; 
    wire core_id_ctrl_decoder_25 ; 
    wire core_id_ctrl_decoder_26 ; 
    wire[31:0] core_id_ctrl_decoder_decoded_plaInput ; 
    wire[31:0] core_id_ctrl_decoder_decoded_invInputs =~ core_id_ctrl_decoder_decoded_plaInput ; 
    wire[39:0] core_id_ctrl_decoder_decoded_invMatrixOutputs ; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_1 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_2 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_3 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_4 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_5 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_6 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_7 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_8 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_9 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_10 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_11 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_12 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_13 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_14 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_15 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_16 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_17 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_18 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_19 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_20 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_21 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_22 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_23 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_24 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_25 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_26 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_27 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_28 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_29 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_30 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_31 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_32 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_33 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_34 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_35 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_36 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_37 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_38 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_39 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_40 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_41 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_42 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_43 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_44 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_45 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_46 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_47 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_48 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_49 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_50 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_51 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_52 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_53 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_54 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_55 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_56 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_57 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_58 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_59 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_60 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_61 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_62 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_64 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_65 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_66 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_67 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_69 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_70 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_1 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_2 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_3 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_4 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_5 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_6 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_7 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_8 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_9 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_10 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_11 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_12 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_13 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_14 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_15 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_16 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_17 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_19 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_20 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_21 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_22 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_23 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_24 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_25 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_26 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_27 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_28 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_29 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_30 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_31 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_32 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_33 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_34 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_35 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_36 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_37 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_38 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_39 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_40 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_41 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_42 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_43 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_44 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_45 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_46 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_47 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_48 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_49 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_50 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_51 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_52 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_53 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_54 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_55 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_56 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_57 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_58 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_60 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_61 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_62 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_64 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_65 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_66 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_67 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_69 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_70 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_1 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_2 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_3 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_4 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_8 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_9 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_10 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_11 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_12 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_13 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_14 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_19 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_21 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_22 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_23 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_24 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_25 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_26 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_27 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_28 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_30 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_31 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_32 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_33 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_34 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_35 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_36 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_37 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_38 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_39 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_40 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_41 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_42 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_43 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_44 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_45 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_46 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_47 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_48 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_49 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_50 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_51 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_52 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_53 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_54 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_55 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_60 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_64 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_65 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_67 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_69 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_1 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_2 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_3 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_4 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_6 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_7 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_8 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_9 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_10 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_11 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_12 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_13 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_14 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_15 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_16 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_19 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_21 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_22 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_23 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_24 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_25 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_26 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_27 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_28 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_30 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_31 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_32 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_33 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_34 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_35 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_36 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_37 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_38 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_39 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_40 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_41 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_42 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_43 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_44 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_45 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_46 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_47 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_48 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_49 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_50 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_51 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_52 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_53 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_54 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_55 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_60 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_64 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_65 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_67 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_69 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_2 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_4 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_5 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_8 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_9 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_10 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_13 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_14 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_15 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_16 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_17 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_20 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_24 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_29 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_38 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_45 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_50 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_56 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_57 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_58 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_61 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_62 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_66 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_70 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_1 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_3 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_5 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_7 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_20 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_22 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_27 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_28 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_34 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_36 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_40 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_47 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_52 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_1 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_2 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_3 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_4 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_5 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_6 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_6 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_7 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_9 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_10 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_11 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_19 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_21 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_21 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_26 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_27 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_28 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_29 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_30 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_33 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_34 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_35 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_36 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_39 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_39 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_41 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_41 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_42 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_46 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_47 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_51 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_52 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_53 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_54 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_55 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_56 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_57 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_60 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_61 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_64 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_65 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_67 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_69 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_1 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_4 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_5 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_8 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_8 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_3 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_11 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_12 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_13 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_7 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_2 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_2 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_10 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_18 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_12 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_20 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_13 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_22 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_36 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_25 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_38 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_27 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_23 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_22 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_30 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_25 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_48 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_64 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_35 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_29 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_6 , core_id_ctrl_decoder_decoded_andMatrixInput_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_4 , core_id_ctrl_decoder_decoded_andMatrixInput_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo ={ core_id_ctrl_decoder_decoded_lo_hi , core_id_ctrl_decoder_decoded_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_2 , core_id_ctrl_decoder_decoded_andMatrixInput_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_0 , core_id_ctrl_decoder_decoded_andMatrixInput_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi ={ core_id_ctrl_decoder_decoded_hi_hi , core_id_ctrl_decoder_decoded_hi_lo }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T ={ core_id_ctrl_decoder_decoded_hi , core_id_ctrl_decoder_decoded_lo }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_1 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_2 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_3 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_6 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_9 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_14 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_14 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_3 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_3 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_26 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_33 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_53 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_55 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_26 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_23 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_58 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_59 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_46 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_27 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_62 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_63 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_51 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_32 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_67 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_1 , core_id_ctrl_decoder_decoded_andMatrixInput_7_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_1 , core_id_ctrl_decoder_decoded_andMatrixInput_5_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_1 ={ core_id_ctrl_decoder_decoded_lo_hi_1 , core_id_ctrl_decoder_decoded_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_1 , core_id_ctrl_decoder_decoded_andMatrixInput_3_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_1 , core_id_ctrl_decoder_decoded_andMatrixInput_1_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_1 ={ core_id_ctrl_decoder_decoded_hi_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_1 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_3 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_4 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_1 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_7 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_6 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_14 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_15 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_8 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_18 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_19 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_23 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_25 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_23 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_19 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_28 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_29 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_27 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_22 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_32 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_33 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_32 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_26 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_37 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_2 , core_id_ctrl_decoder_decoded_andMatrixInput_7_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_2 , core_id_ctrl_decoder_decoded_andMatrixInput_5_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_2 ={ core_id_ctrl_decoder_decoded_lo_hi_2 , core_id_ctrl_decoder_decoded_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_2 , core_id_ctrl_decoder_decoded_andMatrixInput_3_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_2 , core_id_ctrl_decoder_decoded_andMatrixInput_1_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_2 ={ core_id_ctrl_decoder_decoded_hi_hi_2 , core_id_ctrl_decoder_decoded_hi_lo_2 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_4 ={ core_id_ctrl_decoder_decoded_hi_2 , core_id_ctrl_decoder_decoded_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_3 , core_id_ctrl_decoder_decoded_andMatrixInput_7_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_3 , core_id_ctrl_decoder_decoded_andMatrixInput_5_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_3 ={ core_id_ctrl_decoder_decoded_lo_hi_3 , core_id_ctrl_decoder_decoded_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_3 , core_id_ctrl_decoder_decoded_andMatrixInput_3_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_3 , core_id_ctrl_decoder_decoded_andMatrixInput_1_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_3 ={ core_id_ctrl_decoder_decoded_hi_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_3 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_6 ={ core_id_ctrl_decoder_decoded_hi_3 , core_id_ctrl_decoder_decoded_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_4 , core_id_ctrl_decoder_decoded_andMatrixInput_7_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_4 , core_id_ctrl_decoder_decoded_andMatrixInput_5_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_4 ={ core_id_ctrl_decoder_decoded_lo_hi_4 , core_id_ctrl_decoder_decoded_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_4 , core_id_ctrl_decoder_decoded_andMatrixInput_3_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_4 , core_id_ctrl_decoder_decoded_andMatrixInput_1_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_4 ={ core_id_ctrl_decoder_decoded_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_lo_4 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_8 ={ core_id_ctrl_decoder_decoded_hi_4 , core_id_ctrl_decoder_decoded_lo_4 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_5 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_6 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_7 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_16 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_17 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_20 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_29 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_56 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_57 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_58 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_61 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_62 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_66 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_70 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_5 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_17 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_20 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_29 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_56 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_57 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_58 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_61 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_62 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_66 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_70 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_5 , core_id_ctrl_decoder_decoded_andMatrixInput_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_5 , core_id_ctrl_decoder_decoded_andMatrixInput_6_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_5 ={ core_id_ctrl_decoder_decoded_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_5 , core_id_ctrl_decoder_decoded_andMatrixInput_4_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_5 , core_id_ctrl_decoder_decoded_andMatrixInput_1_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_5 ={ core_id_ctrl_decoder_decoded_hi_hi_hi , core_id_ctrl_decoder_decoded_andMatrixInput_2_5 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_5 ={ core_id_ctrl_decoder_decoded_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_5 }; 
    wire[8:0] core__id_ctrl_decoder_decoded_T_10 ={ core_id_ctrl_decoder_decoded_hi_5 , core_id_ctrl_decoder_decoded_lo_5 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_6 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_7 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_11 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_12 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_18 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_19 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_21 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_22 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_26 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_27 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_28 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_30 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_31 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_32 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_33 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_34 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_35 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_36 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_37 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_39 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_40 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_41 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_42 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_43 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_46 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_47 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_48 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_51 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_52 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_53 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_54 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_55 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_59 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_60 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_63 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_64 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_65 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_67 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_68 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_69 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_6 , core_id_ctrl_decoder_decoded_andMatrixInput_4_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_6 ={ core_id_ctrl_decoder_decoded_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_5_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_6 , core_id_ctrl_decoder_decoded_andMatrixInput_1_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_6 ={ core_id_ctrl_decoder_decoded_hi_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_2_6 }; 
    wire[5:0] core__id_ctrl_decoder_decoded_T_12 ={ core_id_ctrl_decoder_decoded_hi_6 , core_id_ctrl_decoder_decoded_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_7 , core_id_ctrl_decoder_decoded_andMatrixInput_5_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_7 ={ core_id_ctrl_decoder_decoded_lo_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_6_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_7 , core_id_ctrl_decoder_decoded_andMatrixInput_3_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_7 , core_id_ctrl_decoder_decoded_andMatrixInput_1_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_7 ={ core_id_ctrl_decoder_decoded_hi_hi_7 , core_id_ctrl_decoder_decoded_hi_lo_6 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_8 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_9 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_10 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_11 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_12 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_13 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_14 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_15 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_16 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_17 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_18 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_19 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_23 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_24 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_25 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_26 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_29 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_30 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_31 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_32 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_33 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_35 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_37 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_38 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_42 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_43 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_44 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_45 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_46 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_48 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_49 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_50 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_51 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_53 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_54 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_55 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_56 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_57 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_58 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_59 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_60 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_61 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_62 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_63 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_64 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_65 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_66 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_68 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_69 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_70 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_6 , core_id_ctrl_decoder_decoded_andMatrixInput_8_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_8 , core_id_ctrl_decoder_decoded_andMatrixInput_6_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_8 ={ core_id_ctrl_decoder_decoded_lo_hi_8 , core_id_ctrl_decoder_decoded_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_8 , core_id_ctrl_decoder_decoded_andMatrixInput_4_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_8 , core_id_ctrl_decoder_decoded_andMatrixInput_1_8 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_8 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_2_8 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_8 ={ core_id_ctrl_decoder_decoded_hi_hi_8 , core_id_ctrl_decoder_decoded_hi_lo_7 }; 
    wire[8:0] core__id_ctrl_decoder_decoded_T_16 ={ core_id_ctrl_decoder_decoded_hi_8 , core_id_ctrl_decoder_decoded_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_8 , core_id_ctrl_decoder_decoded_andMatrixInput_7_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_9 , core_id_ctrl_decoder_decoded_andMatrixInput_5_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_9 ={ core_id_ctrl_decoder_decoded_lo_hi_9 , core_id_ctrl_decoder_decoded_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_9 , core_id_ctrl_decoder_decoded_andMatrixInput_3_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_9 , core_id_ctrl_decoder_decoded_andMatrixInput_1_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_9 ={ core_id_ctrl_decoder_decoded_hi_hi_9 , core_id_ctrl_decoder_decoded_hi_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_8 , core_id_ctrl_decoder_decoded_andMatrixInput_8_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_10 , core_id_ctrl_decoder_decoded_andMatrixInput_6_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_10 ={ core_id_ctrl_decoder_decoded_lo_hi_10 , core_id_ctrl_decoder_decoded_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_10 , core_id_ctrl_decoder_decoded_andMatrixInput_4_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_10 , core_id_ctrl_decoder_decoded_andMatrixInput_1_10 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_10 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_2_10 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_10 ={ core_id_ctrl_decoder_decoded_hi_hi_10 , core_id_ctrl_decoder_decoded_hi_lo_9 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_1 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_11 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_7 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_17 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_10 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_13 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_12 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_15 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_14 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_2 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_3 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_4 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_5 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_29 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_34 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_10 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_1 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_6 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_5 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_9 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_8 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_11 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_23 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_11 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_12 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_13 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_14 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_17 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_18 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_36 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_21 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_22 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_2 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_3 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_4 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_5 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_29 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_31 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_6 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_7 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_4 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_1 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_4 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_5 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_6 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_7 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_8 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_9 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_12 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_11 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_11 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_13 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_13 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_15 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_16 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_20 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_18 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_19 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_20 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_9 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_2 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_3 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_26 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_4 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_5 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_28 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_30 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_31 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_34 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_1 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_1 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_4 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_5 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_6 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_7 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_7 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_9 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_10 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_10 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_10 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_12 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_12 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_15 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_16 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_17 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_18 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_19 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_26 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_26 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_30 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_30 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_34 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_1 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_4 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_4 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_6 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_6 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_8 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_10 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_9 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_9 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_11 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_11 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_14 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_15 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_17 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_17 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_18 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_20 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_16 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_2 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_24 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_23 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_27 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_1 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_3 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_3 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_5 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_4 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_7 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_8 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_8 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_5 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_6 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_7 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_12 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_13 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_15 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_14 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_15 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_18 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30_1 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_20 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_4 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_31 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_8 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_15 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_6 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_31_1 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_14 , core_id_ctrl_decoder_decoded_andMatrixInput_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_12 , core_id_ctrl_decoder_decoded_andMatrixInput_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_9 ={ core_id_ctrl_decoder_decoded_lo_lo_hi , core_id_ctrl_decoder_decoded_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_10 , core_id_ctrl_decoder_decoded_andMatrixInput_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_3 , core_id_ctrl_decoder_decoded_andMatrixInput_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_11 ={ core_id_ctrl_decoder_decoded_lo_hi_hi , core_id_ctrl_decoder_decoded_lo_hi_lo }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_11 ={ core_id_ctrl_decoder_decoded_lo_hi_11 , core_id_ctrl_decoder_decoded_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_10 , core_id_ctrl_decoder_decoded_andMatrixInput_7_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_11 , core_id_ctrl_decoder_decoded_andMatrixInput_5_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_10 ={ core_id_ctrl_decoder_decoded_hi_lo_hi , core_id_ctrl_decoder_decoded_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_11 , core_id_ctrl_decoder_decoded_andMatrixInput_3_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_11 , core_id_ctrl_decoder_decoded_andMatrixInput_1_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_11 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_hi_hi_lo }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_11 ={ core_id_ctrl_decoder_decoded_hi_hi_11 , core_id_ctrl_decoder_decoded_hi_lo_10 }; 
    wire[15:0] core__id_ctrl_decoder_decoded_T_22 ={ core_id_ctrl_decoder_decoded_hi_11 , core_id_ctrl_decoder_decoded_lo_11 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_1 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_3 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_4 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_5 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_6 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_7 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_9 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_10 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_13 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_14 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_16 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_16 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_17 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_19 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_8 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29_1 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_23 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_4 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_1 , core_id_ctrl_decoder_decoded_andMatrixInput_11_1 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_10 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_12_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_10 , core_id_ctrl_decoder_decoded_andMatrixInput_8_4 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_12 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_9_1 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_12 ={ core_id_ctrl_decoder_decoded_lo_hi_12 , core_id_ctrl_decoder_decoded_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_12 , core_id_ctrl_decoder_decoded_andMatrixInput_5_12 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_11 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_6_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_12 , core_id_ctrl_decoder_decoded_andMatrixInput_3_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_12 , core_id_ctrl_decoder_decoded_andMatrixInput_1_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_12 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_hi_lo_1 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_12 ={ core_id_ctrl_decoder_decoded_hi_hi_12 , core_id_ctrl_decoder_decoded_hi_lo_11 }; 
    wire[12:0] core__id_ctrl_decoder_decoded_T_24 ={ core_id_ctrl_decoder_decoded_hi_12 , core_id_ctrl_decoder_decoded_lo_12 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_12 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_13 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_15 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_15 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_16 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_18 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_18 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_23 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_23 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_25 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_25 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_31 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_32 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_37 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_44 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_44 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_45 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_49 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_49 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_50 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_59 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_59 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_63 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_63 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_68 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_68 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_12 , core_id_ctrl_decoder_decoded_andMatrixInput_7_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_13 , core_id_ctrl_decoder_decoded_andMatrixInput_5_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_13 ={ core_id_ctrl_decoder_decoded_lo_hi_13 , core_id_ctrl_decoder_decoded_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_13 , core_id_ctrl_decoder_decoded_andMatrixInput_3_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_13 , core_id_ctrl_decoder_decoded_andMatrixInput_1_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_13 ={ core_id_ctrl_decoder_decoded_hi_hi_13 , core_id_ctrl_decoder_decoded_hi_lo_12 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_26 ={ core_id_ctrl_decoder_decoded_hi_13 , core_id_ctrl_decoder_decoded_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_12 , core_id_ctrl_decoder_decoded_andMatrixInput_8_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_14 , core_id_ctrl_decoder_decoded_andMatrixInput_6_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_14 ={ core_id_ctrl_decoder_decoded_lo_hi_14 , core_id_ctrl_decoder_decoded_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_14 , core_id_ctrl_decoder_decoded_andMatrixInput_4_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_14 , core_id_ctrl_decoder_decoded_andMatrixInput_1_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_14 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_andMatrixInput_2_14 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_14 ={ core_id_ctrl_decoder_decoded_hi_hi_14 , core_id_ctrl_decoder_decoded_hi_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_13 , core_id_ctrl_decoder_decoded_andMatrixInput_8_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_15 , core_id_ctrl_decoder_decoded_andMatrixInput_6_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_15 ={ core_id_ctrl_decoder_decoded_lo_hi_15 , core_id_ctrl_decoder_decoded_lo_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_15 , core_id_ctrl_decoder_decoded_andMatrixInput_4_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_15 , core_id_ctrl_decoder_decoded_andMatrixInput_1_15 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_15 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_2_15 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_15 ={ core_id_ctrl_decoder_decoded_hi_hi_15 , core_id_ctrl_decoder_decoded_hi_lo_14 }; 
    wire[8:0] core__id_ctrl_decoder_decoded_T_30 ={ core_id_ctrl_decoder_decoded_hi_15 , core_id_ctrl_decoder_decoded_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_7 , core_id_ctrl_decoder_decoded_andMatrixInput_9_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_16 , core_id_ctrl_decoder_decoded_andMatrixInput_6_15 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_16 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_7_14 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_16 ={ core_id_ctrl_decoder_decoded_lo_hi_16 , core_id_ctrl_decoder_decoded_lo_lo_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_16 , core_id_ctrl_decoder_decoded_andMatrixInput_4_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_16 , core_id_ctrl_decoder_decoded_andMatrixInput_1_16 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_16 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_2_16 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_16 ={ core_id_ctrl_decoder_decoded_hi_hi_16 , core_id_ctrl_decoder_decoded_hi_lo_15 }; 
    wire[9:0] core__id_ctrl_decoder_decoded_T_32 ={ core_id_ctrl_decoder_decoded_hi_16 , core_id_ctrl_decoder_decoded_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_17 , core_id_ctrl_decoder_decoded_andMatrixInput_5_17 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_17 ={ core_id_ctrl_decoder_decoded_lo_hi_17 , core_id_ctrl_decoder_decoded_andMatrixInput_6_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_17 , core_id_ctrl_decoder_decoded_andMatrixInput_3_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_17 , core_id_ctrl_decoder_decoded_andMatrixInput_1_17 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_17 ={ core_id_ctrl_decoder_decoded_hi_hi_17 , core_id_ctrl_decoder_decoded_hi_lo_16 }; 
    wire[6:0] core__id_ctrl_decoder_decoded_T_34 ={ core_id_ctrl_decoder_decoded_hi_17 , core_id_ctrl_decoder_decoded_lo_17 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_18 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_16 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_59 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_57 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_63 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_61 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_68 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_66 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_18 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_9 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_59 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_43 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_63 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_47 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_68 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_52 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_17 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_4 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_58 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_27 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_63 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_31 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_68 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_36 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_15 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_3 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_56 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_24 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_62 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_28 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_67 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_33 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_8 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_3 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_42 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_24 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_60 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_28 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_65 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_33 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_2 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_2 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_22 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_11 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_27 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_13 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_32 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_17 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_1 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_1 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_21 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_5 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_26 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_7 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_31 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_10 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_1 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_1 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_18 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_4 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_24 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_6 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_28 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_8 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_1 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_1 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_10 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_4 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_21 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_6 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_25 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_8 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_1 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_4 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_4 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_12 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_6 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_16 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_8 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_1 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_40 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_22 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_3 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_3 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_1 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_24 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_21 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_5 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_5 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_7 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_7 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_1 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_21 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_20 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_2 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_3 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_5 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_5 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_7 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_7 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_1 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_21 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_17 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_2 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_3 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_4 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_5 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_25 , core_id_ctrl_decoder_decoded_andMatrixInput_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_1 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_23 , core_id_ctrl_decoder_decoded_andMatrixInput_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_21 , core_id_ctrl_decoder_decoded_andMatrixInput_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_2 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_lo_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_15 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_18 , core_id_ctrl_decoder_decoded_andMatrixInput_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_1 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_16 , core_id_ctrl_decoder_decoded_andMatrixInput_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_1 , core_id_ctrl_decoder_decoded_andMatrixInput_15_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_lo_hi_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_18 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_lo_hi_lo_1 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_18 ={ core_id_ctrl_decoder_decoded_lo_hi_18 , core_id_ctrl_decoder_decoded_lo_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_2 , core_id_ctrl_decoder_decoded_andMatrixInput_12_2 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_1 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_13_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_3 , core_id_ctrl_decoder_decoded_andMatrixInput_10_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_15 , core_id_ctrl_decoder_decoded_andMatrixInput_8_8 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_hi_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_17 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_18 , core_id_ctrl_decoder_decoded_andMatrixInput_5_18 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_6_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_18 , core_id_ctrl_decoder_decoded_andMatrixInput_3_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_18 , core_id_ctrl_decoder_decoded_andMatrixInput_1_18 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_hi_hi_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_18 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_hi_hi_lo_2 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_18 ={ core_id_ctrl_decoder_decoded_hi_hi_18 , core_id_ctrl_decoder_decoded_hi_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28 , core_id_ctrl_decoder_decoded_andMatrixInput_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_2 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_1 , core_id_ctrl_decoder_decoded_andMatrixInput_27_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_1 , core_id_ctrl_decoder_decoded_andMatrixInput_25_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_3 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_1 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_16 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_3 , core_id_ctrl_decoder_decoded_lo_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_1 , core_id_ctrl_decoder_decoded_andMatrixInput_23_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_1 , core_id_ctrl_decoder_decoded_andMatrixInput_21_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_2 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_1 , core_id_ctrl_decoder_decoded_andMatrixInput_19_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_1 , core_id_ctrl_decoder_decoded_andMatrixInput_17_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_1 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_19 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_lo_hi_lo_2 }; 
    wire[14:0] core_id_ctrl_decoder_decoded_lo_19 ={ core_id_ctrl_decoder_decoded_lo_hi_19 , core_id_ctrl_decoder_decoded_lo_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_2 , core_id_ctrl_decoder_decoded_andMatrixInput_15_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_3 , core_id_ctrl_decoder_decoded_andMatrixInput_13_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_2 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_3 , core_id_ctrl_decoder_decoded_andMatrixInput_11_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_9 , core_id_ctrl_decoder_decoded_andMatrixInput_9_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_3 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_18 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_18 , core_id_ctrl_decoder_decoded_andMatrixInput_7_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_19 , core_id_ctrl_decoder_decoded_andMatrixInput_5_19 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_3 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_19 , core_id_ctrl_decoder_decoded_andMatrixInput_3_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_19 , core_id_ctrl_decoder_decoded_andMatrixInput_1_19 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_9 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_1 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_19 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_9 , core_id_ctrl_decoder_decoded_hi_hi_lo_3 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_19 ={ core_id_ctrl_decoder_decoded_hi_hi_19 , core_id_ctrl_decoder_decoded_hi_lo_18 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_17 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_20 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_19 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_22 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_21 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_24 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_23 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_31 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_32 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_38 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_37 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_40 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_39 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_40 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_43 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_42 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_43 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_49 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_51 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_66 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_10 , core_id_ctrl_decoder_decoded_andMatrixInput_9_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_20 , core_id_ctrl_decoder_decoded_andMatrixInput_6_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_20 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_andMatrixInput_7_17 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_20 ={ core_id_ctrl_decoder_decoded_lo_hi_20 , core_id_ctrl_decoder_decoded_lo_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_20 , core_id_ctrl_decoder_decoded_andMatrixInput_4_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_20 , core_id_ctrl_decoder_decoded_andMatrixInput_1_20 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_20 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_10 , core_id_ctrl_decoder_decoded_andMatrixInput_2_20 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_20 ={ core_id_ctrl_decoder_decoded_hi_hi_20 , core_id_ctrl_decoder_decoded_hi_lo_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_4 , core_id_ctrl_decoder_decoded_andMatrixInput_13_3 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_18 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_14_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_4 , core_id_ctrl_decoder_decoded_andMatrixInput_11_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_11 , core_id_ctrl_decoder_decoded_andMatrixInput_9_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_21 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_lo_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_21 ={ core_id_ctrl_decoder_decoded_lo_hi_21 , core_id_ctrl_decoder_decoded_lo_lo_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_20 , core_id_ctrl_decoder_decoded_andMatrixInput_7_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_21 , core_id_ctrl_decoder_decoded_andMatrixInput_5_21 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_20 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_21 , core_id_ctrl_decoder_decoded_andMatrixInput_3_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_21 , core_id_ctrl_decoder_decoded_andMatrixInput_1_21 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_21 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_11 , core_id_ctrl_decoder_decoded_hi_hi_lo_4 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_21 ={ core_id_ctrl_decoder_decoded_hi_hi_21 , core_id_ctrl_decoder_decoded_hi_lo_20 }; 
    wire[14:0] core__id_ctrl_decoder_decoded_T_42 ={ core_id_ctrl_decoder_decoded_hi_21 , core_id_ctrl_decoder_decoded_lo_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_4 , core_id_ctrl_decoder_decoded_andMatrixInput_15_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_5 , core_id_ctrl_decoder_decoded_andMatrixInput_13_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_19 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_5 , core_id_ctrl_decoder_decoded_andMatrixInput_11_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_12 , core_id_ctrl_decoder_decoded_andMatrixInput_9_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_22 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_lo_hi_lo_4 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_22 ={ core_id_ctrl_decoder_decoded_lo_hi_22 , core_id_ctrl_decoder_decoded_lo_lo_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_21 , core_id_ctrl_decoder_decoded_andMatrixInput_7_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_22 , core_id_ctrl_decoder_decoded_andMatrixInput_5_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_21 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_22 , core_id_ctrl_decoder_decoded_andMatrixInput_3_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_22 , core_id_ctrl_decoder_decoded_andMatrixInput_1_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_22 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_12 , core_id_ctrl_decoder_decoded_hi_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_22 ={ core_id_ctrl_decoder_decoded_hi_hi_22 , core_id_ctrl_decoder_decoded_hi_lo_21 }; 
    wire[15:0] core__id_ctrl_decoder_decoded_T_44 ={ core_id_ctrl_decoder_decoded_hi_22 , core_id_ctrl_decoder_decoded_lo_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_22 , core_id_ctrl_decoder_decoded_andMatrixInput_7_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_23 , core_id_ctrl_decoder_decoded_andMatrixInput_5_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_23 ={ core_id_ctrl_decoder_decoded_lo_hi_23 , core_id_ctrl_decoder_decoded_lo_lo_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_23 , core_id_ctrl_decoder_decoded_andMatrixInput_3_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_23 , core_id_ctrl_decoder_decoded_andMatrixInput_1_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_23 ={ core_id_ctrl_decoder_decoded_hi_hi_23 , core_id_ctrl_decoder_decoded_hi_lo_22 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_46 ={ core_id_ctrl_decoder_decoded_hi_23 , core_id_ctrl_decoder_decoded_lo_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_21 , core_id_ctrl_decoder_decoded_andMatrixInput_8_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_24 , core_id_ctrl_decoder_decoded_andMatrixInput_6_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_24 ={ core_id_ctrl_decoder_decoded_lo_hi_24 , core_id_ctrl_decoder_decoded_lo_lo_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_24 , core_id_ctrl_decoder_decoded_andMatrixInput_4_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_24 , core_id_ctrl_decoder_decoded_andMatrixInput_1_24 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_24 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_13 , core_id_ctrl_decoder_decoded_andMatrixInput_2_24 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_24 ={ core_id_ctrl_decoder_decoded_hi_hi_24 , core_id_ctrl_decoder_decoded_hi_lo_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_22 , core_id_ctrl_decoder_decoded_andMatrixInput_8_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_25 , core_id_ctrl_decoder_decoded_andMatrixInput_6_24 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_25 ={ core_id_ctrl_decoder_decoded_lo_hi_25 , core_id_ctrl_decoder_decoded_lo_lo_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_25 , core_id_ctrl_decoder_decoded_andMatrixInput_4_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_25 , core_id_ctrl_decoder_decoded_andMatrixInput_1_25 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_25 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_14 , core_id_ctrl_decoder_decoded_andMatrixInput_2_25 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_25 ={ core_id_ctrl_decoder_decoded_hi_hi_25 , core_id_ctrl_decoder_decoded_hi_lo_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_25 , core_id_ctrl_decoder_decoded_andMatrixInput_7_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_26 , core_id_ctrl_decoder_decoded_andMatrixInput_5_26 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_26 ={ core_id_ctrl_decoder_decoded_lo_hi_26 , core_id_ctrl_decoder_decoded_lo_lo_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_26 , core_id_ctrl_decoder_decoded_andMatrixInput_3_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_26 , core_id_ctrl_decoder_decoded_andMatrixInput_1_26 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_26 ={ core_id_ctrl_decoder_decoded_hi_hi_26 , core_id_ctrl_decoder_decoded_hi_lo_25 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_52 ={ core_id_ctrl_decoder_decoded_hi_26 , core_id_ctrl_decoder_decoded_lo_26 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_24 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_25 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_16 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_27 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_28 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_29 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_30 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_20 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_21 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_44 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_45 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_48 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_47 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_48 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_35 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_52 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_39 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_41 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_44 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_45 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_49 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_53 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_26 , core_id_ctrl_decoder_decoded_andMatrixInput_7_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_27 , core_id_ctrl_decoder_decoded_andMatrixInput_5_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_27 ={ core_id_ctrl_decoder_decoded_lo_hi_27 , core_id_ctrl_decoder_decoded_lo_lo_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_27 , core_id_ctrl_decoder_decoded_andMatrixInput_3_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_27 , core_id_ctrl_decoder_decoded_andMatrixInput_1_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_27 ={ core_id_ctrl_decoder_decoded_hi_hi_27 , core_id_ctrl_decoder_decoded_hi_lo_26 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_54 ={ core_id_ctrl_decoder_decoded_hi_27 , core_id_ctrl_decoder_decoded_lo_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_25 , core_id_ctrl_decoder_decoded_andMatrixInput_8_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_28 , core_id_ctrl_decoder_decoded_andMatrixInput_6_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_28 ={ core_id_ctrl_decoder_decoded_lo_hi_28 , core_id_ctrl_decoder_decoded_lo_lo_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_28 , core_id_ctrl_decoder_decoded_andMatrixInput_4_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_28 , core_id_ctrl_decoder_decoded_andMatrixInput_1_28 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_28 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_15 , core_id_ctrl_decoder_decoded_andMatrixInput_2_28 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_28 ={ core_id_ctrl_decoder_decoded_hi_hi_28 , core_id_ctrl_decoder_decoded_hi_lo_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_8 , core_id_ctrl_decoder_decoded_andMatrixInput_10_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_26 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_11_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_28 , core_id_ctrl_decoder_decoded_andMatrixInput_7_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_29 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_8 , core_id_ctrl_decoder_decoded_andMatrixInput_8_16 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_29 ={ core_id_ctrl_decoder_decoded_lo_hi_29 , core_id_ctrl_decoder_decoded_lo_lo_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_29 , core_id_ctrl_decoder_decoded_andMatrixInput_4_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_28 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_5_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_29 , core_id_ctrl_decoder_decoded_andMatrixInput_1_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_29 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_16 , core_id_ctrl_decoder_decoded_andMatrixInput_2_29 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_hi_29 ={ core_id_ctrl_decoder_decoded_hi_hi_29 , core_id_ctrl_decoder_decoded_hi_lo_28 }; 
    wire[11:0] core__id_ctrl_decoder_decoded_T_58 ={ core_id_ctrl_decoder_decoded_hi_29 , core_id_ctrl_decoder_decoded_lo_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_6 , core_id_ctrl_decoder_decoded_andMatrixInput_13_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_27 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_14_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_7 , core_id_ctrl_decoder_decoded_andMatrixInput_11_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_17 , core_id_ctrl_decoder_decoded_andMatrixInput_9_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_30 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_9 , core_id_ctrl_decoder_decoded_lo_hi_lo_5 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_30 ={ core_id_ctrl_decoder_decoded_lo_hi_30 , core_id_ctrl_decoder_decoded_lo_lo_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_29 , core_id_ctrl_decoder_decoded_andMatrixInput_7_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_30 , core_id_ctrl_decoder_decoded_andMatrixInput_5_30 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_29 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_hi_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_30 , core_id_ctrl_decoder_decoded_andMatrixInput_3_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_30 , core_id_ctrl_decoder_decoded_andMatrixInput_1_30 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_30 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_17 , core_id_ctrl_decoder_decoded_hi_hi_lo_6 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_30 ={ core_id_ctrl_decoder_decoded_hi_hi_30 , core_id_ctrl_decoder_decoded_hi_lo_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_6 , core_id_ctrl_decoder_decoded_andMatrixInput_15_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_7 , core_id_ctrl_decoder_decoded_andMatrixInput_13_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_28 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_8 , core_id_ctrl_decoder_decoded_lo_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_8 , core_id_ctrl_decoder_decoded_andMatrixInput_11_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_18 , core_id_ctrl_decoder_decoded_andMatrixInput_9_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_31 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_10 , core_id_ctrl_decoder_decoded_lo_hi_lo_6 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_31 ={ core_id_ctrl_decoder_decoded_lo_hi_31 , core_id_ctrl_decoder_decoded_lo_lo_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_30 , core_id_ctrl_decoder_decoded_andMatrixInput_7_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_31 , core_id_ctrl_decoder_decoded_andMatrixInput_5_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_30 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_8 , core_id_ctrl_decoder_decoded_hi_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_31 , core_id_ctrl_decoder_decoded_andMatrixInput_3_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_31 , core_id_ctrl_decoder_decoded_andMatrixInput_1_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_31 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_18 , core_id_ctrl_decoder_decoded_hi_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_31 ={ core_id_ctrl_decoder_decoded_hi_hi_31 , core_id_ctrl_decoder_decoded_hi_lo_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_31 , core_id_ctrl_decoder_decoded_andMatrixInput_7_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_32 , core_id_ctrl_decoder_decoded_andMatrixInput_5_32 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_32 ={ core_id_ctrl_decoder_decoded_lo_hi_32 , core_id_ctrl_decoder_decoded_lo_lo_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_32 , core_id_ctrl_decoder_decoded_andMatrixInput_3_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_32 , core_id_ctrl_decoder_decoded_andMatrixInput_1_32 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_32 ={ core_id_ctrl_decoder_decoded_hi_hi_32 , core_id_ctrl_decoder_decoded_hi_lo_31 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_64 ={ core_id_ctrl_decoder_decoded_hi_32 , core_id_ctrl_decoder_decoded_lo_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_30 , core_id_ctrl_decoder_decoded_andMatrixInput_8_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_33 , core_id_ctrl_decoder_decoded_andMatrixInput_6_32 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_33 ={ core_id_ctrl_decoder_decoded_lo_hi_33 , core_id_ctrl_decoder_decoded_lo_lo_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_33 , core_id_ctrl_decoder_decoded_andMatrixInput_4_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_33 , core_id_ctrl_decoder_decoded_andMatrixInput_1_33 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_33 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_19 , core_id_ctrl_decoder_decoded_andMatrixInput_2_33 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_33 ={ core_id_ctrl_decoder_decoded_hi_hi_33 , core_id_ctrl_decoder_decoded_hi_lo_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_31 , core_id_ctrl_decoder_decoded_andMatrixInput_8_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_34 , core_id_ctrl_decoder_decoded_andMatrixInput_6_33 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_34 ={ core_id_ctrl_decoder_decoded_lo_hi_34 , core_id_ctrl_decoder_decoded_lo_lo_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_34 , core_id_ctrl_decoder_decoded_andMatrixInput_4_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_34 , core_id_ctrl_decoder_decoded_andMatrixInput_1_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_34 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_20 , core_id_ctrl_decoder_decoded_andMatrixInput_2_34 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_34 ={ core_id_ctrl_decoder_decoded_hi_hi_34 , core_id_ctrl_decoder_decoded_hi_lo_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_8 , core_id_ctrl_decoder_decoded_andMatrixInput_13_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_32 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_9 , core_id_ctrl_decoder_decoded_andMatrixInput_14_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_9 , core_id_ctrl_decoder_decoded_andMatrixInput_11_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_21 , core_id_ctrl_decoder_decoded_andMatrixInput_9_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_35 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_11 , core_id_ctrl_decoder_decoded_lo_hi_lo_7 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_35 ={ core_id_ctrl_decoder_decoded_lo_hi_35 , core_id_ctrl_decoder_decoded_lo_lo_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_34 , core_id_ctrl_decoder_decoded_andMatrixInput_7_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_35 , core_id_ctrl_decoder_decoded_andMatrixInput_5_35 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_34 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_9 , core_id_ctrl_decoder_decoded_hi_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_35 , core_id_ctrl_decoder_decoded_andMatrixInput_3_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_35 , core_id_ctrl_decoder_decoded_andMatrixInput_1_35 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_35 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_21 , core_id_ctrl_decoder_decoded_hi_hi_lo_8 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_35 ={ core_id_ctrl_decoder_decoded_hi_hi_35 , core_id_ctrl_decoder_decoded_hi_lo_34 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_22 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_34 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_35 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_24 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_14 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_26 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_16 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_28 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_41 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_29 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_30 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_31 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_32 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_46 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_33 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_34 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_19 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_50 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_33 , core_id_ctrl_decoder_decoded_andMatrixInput_8_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_36 , core_id_ctrl_decoder_decoded_andMatrixInput_6_35 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_36 ={ core_id_ctrl_decoder_decoded_lo_hi_36 , core_id_ctrl_decoder_decoded_lo_lo_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_35 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_36 , core_id_ctrl_decoder_decoded_andMatrixInput_4_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_36 , core_id_ctrl_decoder_decoded_andMatrixInput_1_36 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_36 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_22 , core_id_ctrl_decoder_decoded_andMatrixInput_2_36 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_36 ={ core_id_ctrl_decoder_decoded_hi_hi_36 , core_id_ctrl_decoder_decoded_hi_lo_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_10 , core_id_ctrl_decoder_decoded_andMatrixInput_12_9 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_34 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_10 , core_id_ctrl_decoder_decoded_andMatrixInput_13_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_12 , core_id_ctrl_decoder_decoded_andMatrixInput_10_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_34 , core_id_ctrl_decoder_decoded_andMatrixInput_8_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_37 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_12 , core_id_ctrl_decoder_decoded_lo_hi_lo_8 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_37 ={ core_id_ctrl_decoder_decoded_lo_hi_37 , core_id_ctrl_decoder_decoded_lo_lo_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_37 , core_id_ctrl_decoder_decoded_andMatrixInput_5_37 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_36 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_10 , core_id_ctrl_decoder_decoded_andMatrixInput_6_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_37 , core_id_ctrl_decoder_decoded_andMatrixInput_3_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_37 , core_id_ctrl_decoder_decoded_andMatrixInput_1_37 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_37 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_23 , core_id_ctrl_decoder_decoded_hi_hi_lo_9 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_37 ={ core_id_ctrl_decoder_decoded_hi_hi_37 , core_id_ctrl_decoder_decoded_hi_lo_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_35 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_37 , core_id_ctrl_decoder_decoded_andMatrixInput_7_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_38 , core_id_ctrl_decoder_decoded_andMatrixInput_5_38 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_38 ={ core_id_ctrl_decoder_decoded_lo_hi_38 , core_id_ctrl_decoder_decoded_lo_lo_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_38 , core_id_ctrl_decoder_decoded_andMatrixInput_3_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_38 , core_id_ctrl_decoder_decoded_andMatrixInput_1_38 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_38 ={ core_id_ctrl_decoder_decoded_hi_hi_38 , core_id_ctrl_decoder_decoded_hi_lo_37 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_76 ={ core_id_ctrl_decoder_decoded_hi_38 , core_id_ctrl_decoder_decoded_lo_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_10 , core_id_ctrl_decoder_decoded_andMatrixInput_13_9 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_36 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_11 , core_id_ctrl_decoder_decoded_andMatrixInput_14_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_11 , core_id_ctrl_decoder_decoded_andMatrixInput_11_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_24 , core_id_ctrl_decoder_decoded_andMatrixInput_9_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_39 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_13 , core_id_ctrl_decoder_decoded_lo_hi_lo_9 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_39 ={ core_id_ctrl_decoder_decoded_lo_hi_39 , core_id_ctrl_decoder_decoded_lo_lo_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_38 , core_id_ctrl_decoder_decoded_andMatrixInput_7_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_39 , core_id_ctrl_decoder_decoded_andMatrixInput_5_39 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_38 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_11 , core_id_ctrl_decoder_decoded_hi_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_39 , core_id_ctrl_decoder_decoded_andMatrixInput_3_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_39 , core_id_ctrl_decoder_decoded_andMatrixInput_1_39 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_39 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_24 , core_id_ctrl_decoder_decoded_hi_hi_lo_10 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_39 ={ core_id_ctrl_decoder_decoded_hi_hi_39 , core_id_ctrl_decoder_decoded_hi_lo_38 }; 
    wire[14:0] core__id_ctrl_decoder_decoded_T_78 ={ core_id_ctrl_decoder_decoded_hi_39 , core_id_ctrl_decoder_decoded_lo_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_9 , core_id_ctrl_decoder_decoded_andMatrixInput_15_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_11 , core_id_ctrl_decoder_decoded_andMatrixInput_13_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_37 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_12 , core_id_ctrl_decoder_decoded_lo_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_12 , core_id_ctrl_decoder_decoded_andMatrixInput_11_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_25 , core_id_ctrl_decoder_decoded_andMatrixInput_9_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_40 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_14 , core_id_ctrl_decoder_decoded_lo_hi_lo_10 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_40 ={ core_id_ctrl_decoder_decoded_lo_hi_40 , core_id_ctrl_decoder_decoded_lo_lo_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_39 , core_id_ctrl_decoder_decoded_andMatrixInput_7_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_40 , core_id_ctrl_decoder_decoded_andMatrixInput_5_40 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_39 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_12 , core_id_ctrl_decoder_decoded_hi_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_40 , core_id_ctrl_decoder_decoded_andMatrixInput_3_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_40 , core_id_ctrl_decoder_decoded_andMatrixInput_1_40 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_40 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_25 , core_id_ctrl_decoder_decoded_hi_hi_lo_11 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_40 ={ core_id_ctrl_decoder_decoded_hi_hi_40 , core_id_ctrl_decoder_decoded_hi_lo_39 }; 
    wire[15:0] core__id_ctrl_decoder_decoded_T_80 ={ core_id_ctrl_decoder_decoded_hi_40 , core_id_ctrl_decoder_decoded_lo_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_10 , core_id_ctrl_decoder_decoded_andMatrixInput_15_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_12 , core_id_ctrl_decoder_decoded_andMatrixInput_13_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_38 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_13 , core_id_ctrl_decoder_decoded_lo_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_13 , core_id_ctrl_decoder_decoded_andMatrixInput_11_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_26 , core_id_ctrl_decoder_decoded_andMatrixInput_9_15 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_41 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_15 , core_id_ctrl_decoder_decoded_lo_hi_lo_11 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_41 ={ core_id_ctrl_decoder_decoded_lo_hi_41 , core_id_ctrl_decoder_decoded_lo_lo_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_40 , core_id_ctrl_decoder_decoded_andMatrixInput_7_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_41 , core_id_ctrl_decoder_decoded_andMatrixInput_5_41 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_40 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_13 , core_id_ctrl_decoder_decoded_hi_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_41 , core_id_ctrl_decoder_decoded_andMatrixInput_3_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_41 , core_id_ctrl_decoder_decoded_andMatrixInput_1_41 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_41 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_26 , core_id_ctrl_decoder_decoded_hi_hi_lo_12 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_41 ={ core_id_ctrl_decoder_decoded_hi_hi_41 , core_id_ctrl_decoder_decoded_hi_lo_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_11 , core_id_ctrl_decoder_decoded_andMatrixInput_15_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_13 , core_id_ctrl_decoder_decoded_andMatrixInput_13_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_39 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_14 , core_id_ctrl_decoder_decoded_lo_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_14 , core_id_ctrl_decoder_decoded_andMatrixInput_11_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_27 , core_id_ctrl_decoder_decoded_andMatrixInput_9_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_42 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_16 , core_id_ctrl_decoder_decoded_lo_hi_lo_12 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_42 ={ core_id_ctrl_decoder_decoded_lo_hi_42 , core_id_ctrl_decoder_decoded_lo_lo_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_41 , core_id_ctrl_decoder_decoded_andMatrixInput_7_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_42 , core_id_ctrl_decoder_decoded_andMatrixInput_5_42 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_41 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_14 , core_id_ctrl_decoder_decoded_hi_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_42 , core_id_ctrl_decoder_decoded_andMatrixInput_3_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_42 , core_id_ctrl_decoder_decoded_andMatrixInput_1_42 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_42 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_27 , core_id_ctrl_decoder_decoded_hi_hi_lo_13 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_42 ={ core_id_ctrl_decoder_decoded_hi_hi_42 , core_id_ctrl_decoder_decoded_hi_lo_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_14 , core_id_ctrl_decoder_decoded_andMatrixInput_13_13 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_40 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_15 , core_id_ctrl_decoder_decoded_andMatrixInput_14_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_15 , core_id_ctrl_decoder_decoded_andMatrixInput_11_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_28 , core_id_ctrl_decoder_decoded_andMatrixInput_9_17 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_43 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_17 , core_id_ctrl_decoder_decoded_lo_hi_lo_13 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_43 ={ core_id_ctrl_decoder_decoded_lo_hi_43 , core_id_ctrl_decoder_decoded_lo_lo_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_42 , core_id_ctrl_decoder_decoded_andMatrixInput_7_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_43 , core_id_ctrl_decoder_decoded_andMatrixInput_5_43 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_42 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_15 , core_id_ctrl_decoder_decoded_hi_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_43 , core_id_ctrl_decoder_decoded_andMatrixInput_3_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_43 , core_id_ctrl_decoder_decoded_andMatrixInput_1_43 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_43 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_28 , core_id_ctrl_decoder_decoded_hi_hi_lo_14 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_43 ={ core_id_ctrl_decoder_decoded_hi_hi_43 , core_id_ctrl_decoder_decoded_hi_lo_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_43 , core_id_ctrl_decoder_decoded_andMatrixInput_7_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_44 , core_id_ctrl_decoder_decoded_andMatrixInput_5_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_44 ={ core_id_ctrl_decoder_decoded_lo_hi_44 , core_id_ctrl_decoder_decoded_lo_lo_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_44 , core_id_ctrl_decoder_decoded_andMatrixInput_3_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_44 , core_id_ctrl_decoder_decoded_andMatrixInput_1_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_44 ={ core_id_ctrl_decoder_decoded_hi_hi_44 , core_id_ctrl_decoder_decoded_hi_lo_43 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_88 ={ core_id_ctrl_decoder_decoded_hi_44 , core_id_ctrl_decoder_decoded_lo_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_42 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_42 , core_id_ctrl_decoder_decoded_andMatrixInput_8_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_45 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_45 , core_id_ctrl_decoder_decoded_andMatrixInput_6_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_45 ={ core_id_ctrl_decoder_decoded_lo_hi_45 , core_id_ctrl_decoder_decoded_lo_lo_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_45 , core_id_ctrl_decoder_decoded_andMatrixInput_4_45 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_45 , core_id_ctrl_decoder_decoded_andMatrixInput_1_45 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_45 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_29 , core_id_ctrl_decoder_decoded_andMatrixInput_2_45 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_45 ={ core_id_ctrl_decoder_decoded_hi_hi_45 , core_id_ctrl_decoder_decoded_hi_lo_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_43 , core_id_ctrl_decoder_decoded_andMatrixInput_8_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_46 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_46 , core_id_ctrl_decoder_decoded_andMatrixInput_6_45 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_46 ={ core_id_ctrl_decoder_decoded_lo_hi_46 , core_id_ctrl_decoder_decoded_lo_lo_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_45 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_46 , core_id_ctrl_decoder_decoded_andMatrixInput_4_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_46 , core_id_ctrl_decoder_decoded_andMatrixInput_1_46 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_46 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_30 , core_id_ctrl_decoder_decoded_andMatrixInput_2_46 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_46 ={ core_id_ctrl_decoder_decoded_hi_hi_46 , core_id_ctrl_decoder_decoded_hi_lo_45 }; 
    wire[8:0] core__id_ctrl_decoder_decoded_T_92 ={ core_id_ctrl_decoder_decoded_hi_46 , core_id_ctrl_decoder_decoded_lo_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_44 , core_id_ctrl_decoder_decoded_andMatrixInput_8_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_47 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_47 , core_id_ctrl_decoder_decoded_andMatrixInput_6_46 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_47 ={ core_id_ctrl_decoder_decoded_lo_hi_47 , core_id_ctrl_decoder_decoded_lo_lo_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_46 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_47 , core_id_ctrl_decoder_decoded_andMatrixInput_4_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_47 , core_id_ctrl_decoder_decoded_andMatrixInput_1_47 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_47 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_31 , core_id_ctrl_decoder_decoded_andMatrixInput_2_47 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_47 ={ core_id_ctrl_decoder_decoded_hi_hi_47 , core_id_ctrl_decoder_decoded_hi_lo_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_15 , core_id_ctrl_decoder_decoded_andMatrixInput_13_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_45 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_16 , core_id_ctrl_decoder_decoded_andMatrixInput_14_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_16 , core_id_ctrl_decoder_decoded_andMatrixInput_11_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_32 , core_id_ctrl_decoder_decoded_andMatrixInput_9_18 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_48 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_18 , core_id_ctrl_decoder_decoded_lo_hi_lo_14 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_48 ={ core_id_ctrl_decoder_decoded_lo_hi_48 , core_id_ctrl_decoder_decoded_lo_lo_45 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_47 , core_id_ctrl_decoder_decoded_andMatrixInput_7_45 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_48 , core_id_ctrl_decoder_decoded_andMatrixInput_5_48 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_47 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_16 , core_id_ctrl_decoder_decoded_hi_lo_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_48 , core_id_ctrl_decoder_decoded_andMatrixInput_3_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_48 , core_id_ctrl_decoder_decoded_andMatrixInput_1_48 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_48 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_32 , core_id_ctrl_decoder_decoded_hi_hi_lo_15 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_48 ={ core_id_ctrl_decoder_decoded_hi_hi_48 , core_id_ctrl_decoder_decoded_hi_lo_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_46 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_48 , core_id_ctrl_decoder_decoded_andMatrixInput_7_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_49 , core_id_ctrl_decoder_decoded_andMatrixInput_5_49 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_49 ={ core_id_ctrl_decoder_decoded_lo_hi_49 , core_id_ctrl_decoder_decoded_lo_lo_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_48 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_49 , core_id_ctrl_decoder_decoded_andMatrixInput_3_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_49 , core_id_ctrl_decoder_decoded_andMatrixInput_1_49 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_49 ={ core_id_ctrl_decoder_decoded_hi_hi_49 , core_id_ctrl_decoder_decoded_hi_lo_48 }; 
    wire[7:0] core__id_ctrl_decoder_decoded_T_98 ={ core_id_ctrl_decoder_decoded_hi_49 , core_id_ctrl_decoder_decoded_lo_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_47 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_47 , core_id_ctrl_decoder_decoded_andMatrixInput_8_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_50 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_50 , core_id_ctrl_decoder_decoded_andMatrixInput_6_49 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_50 ={ core_id_ctrl_decoder_decoded_lo_hi_50 , core_id_ctrl_decoder_decoded_lo_lo_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_50 , core_id_ctrl_decoder_decoded_andMatrixInput_4_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_50 , core_id_ctrl_decoder_decoded_andMatrixInput_1_50 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_50 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_33 , core_id_ctrl_decoder_decoded_andMatrixInput_2_50 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_50 ={ core_id_ctrl_decoder_decoded_hi_hi_50 , core_id_ctrl_decoder_decoded_hi_lo_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_48 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_48 , core_id_ctrl_decoder_decoded_andMatrixInput_8_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_51 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_51 , core_id_ctrl_decoder_decoded_andMatrixInput_6_50 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_51 ={ core_id_ctrl_decoder_decoded_lo_hi_51 , core_id_ctrl_decoder_decoded_lo_lo_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_50 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_51 , core_id_ctrl_decoder_decoded_andMatrixInput_4_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_51 , core_id_ctrl_decoder_decoded_andMatrixInput_1_51 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_51 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_34 , core_id_ctrl_decoder_decoded_andMatrixInput_2_51 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_51 ={ core_id_ctrl_decoder_decoded_hi_hi_51 , core_id_ctrl_decoder_decoded_hi_lo_50 }; 
    wire[8:0] core__id_ctrl_decoder_decoded_T_102 ={ core_id_ctrl_decoder_decoded_hi_51 , core_id_ctrl_decoder_decoded_lo_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_35 , core_id_ctrl_decoder_decoded_andMatrixInput_9_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_52 , core_id_ctrl_decoder_decoded_andMatrixInput_6_51 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_52 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_19 , core_id_ctrl_decoder_decoded_andMatrixInput_7_49 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_52 ={ core_id_ctrl_decoder_decoded_lo_hi_52 , core_id_ctrl_decoder_decoded_lo_lo_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_51 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_52 , core_id_ctrl_decoder_decoded_andMatrixInput_4_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_35 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_52 , core_id_ctrl_decoder_decoded_andMatrixInput_1_52 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_52 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_35 , core_id_ctrl_decoder_decoded_andMatrixInput_2_52 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_52 ={ core_id_ctrl_decoder_decoded_hi_hi_52 , core_id_ctrl_decoder_decoded_hi_lo_51 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_50 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_37 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_38 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_6 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_7 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_17 , core_id_ctrl_decoder_decoded_andMatrixInput_12_16 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_50 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_17 , core_id_ctrl_decoder_decoded_andMatrixInput_13_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_20 , core_id_ctrl_decoder_decoded_andMatrixInput_10_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_50 , core_id_ctrl_decoder_decoded_andMatrixInput_8_36 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_53 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_20 , core_id_ctrl_decoder_decoded_lo_hi_lo_15 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_53 ={ core_id_ctrl_decoder_decoded_lo_hi_53 , core_id_ctrl_decoder_decoded_lo_lo_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_53 , core_id_ctrl_decoder_decoded_andMatrixInput_5_53 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_52 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_17 , core_id_ctrl_decoder_decoded_andMatrixInput_6_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_53 , core_id_ctrl_decoder_decoded_andMatrixInput_3_53 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_53 , core_id_ctrl_decoder_decoded_andMatrixInput_1_53 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_53 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_36 , core_id_ctrl_decoder_decoded_hi_hi_lo_16 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_53 ={ core_id_ctrl_decoder_decoded_hi_hi_53 , core_id_ctrl_decoder_decoded_hi_lo_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_17 , core_id_ctrl_decoder_decoded_andMatrixInput_13_16 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_51 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_18 , core_id_ctrl_decoder_decoded_andMatrixInput_14_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_18 , core_id_ctrl_decoder_decoded_andMatrixInput_11_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_37 , core_id_ctrl_decoder_decoded_andMatrixInput_9_21 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_54 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_21 , core_id_ctrl_decoder_decoded_lo_hi_lo_16 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_54 ={ core_id_ctrl_decoder_decoded_lo_hi_54 , core_id_ctrl_decoder_decoded_lo_lo_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_53 , core_id_ctrl_decoder_decoded_andMatrixInput_7_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_54 , core_id_ctrl_decoder_decoded_andMatrixInput_5_54 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_53 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_18 , core_id_ctrl_decoder_decoded_hi_lo_lo_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_54 , core_id_ctrl_decoder_decoded_andMatrixInput_3_54 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_54 , core_id_ctrl_decoder_decoded_andMatrixInput_1_54 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_54 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_37 , core_id_ctrl_decoder_decoded_hi_hi_lo_17 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_54 ={ core_id_ctrl_decoder_decoded_hi_hi_54 , core_id_ctrl_decoder_decoded_hi_lo_53 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_18 , core_id_ctrl_decoder_decoded_andMatrixInput_13_17 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_52 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_19 , core_id_ctrl_decoder_decoded_andMatrixInput_14_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_19 , core_id_ctrl_decoder_decoded_andMatrixInput_11_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_38 , core_id_ctrl_decoder_decoded_andMatrixInput_9_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_55 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_22 , core_id_ctrl_decoder_decoded_lo_hi_lo_17 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_55 ={ core_id_ctrl_decoder_decoded_lo_hi_55 , core_id_ctrl_decoder_decoded_lo_lo_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_54 , core_id_ctrl_decoder_decoded_andMatrixInput_7_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_55 , core_id_ctrl_decoder_decoded_andMatrixInput_5_55 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_54 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_19 , core_id_ctrl_decoder_decoded_hi_lo_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_55 , core_id_ctrl_decoder_decoded_andMatrixInput_3_55 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_55 , core_id_ctrl_decoder_decoded_andMatrixInput_1_55 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_55 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_38 , core_id_ctrl_decoder_decoded_hi_hi_lo_18 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_55 ={ core_id_ctrl_decoder_decoded_hi_hi_55 , core_id_ctrl_decoder_decoded_hi_lo_54 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_20 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_25 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_6 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_7 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_20 , core_id_ctrl_decoder_decoded_andMatrixInput_12_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_53 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_20 , core_id_ctrl_decoder_decoded_andMatrixInput_13_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_23 , core_id_ctrl_decoder_decoded_andMatrixInput_10_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_53 , core_id_ctrl_decoder_decoded_andMatrixInput_8_39 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_56 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_23 , core_id_ctrl_decoder_decoded_lo_hi_lo_18 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_56 ={ core_id_ctrl_decoder_decoded_lo_hi_56 , core_id_ctrl_decoder_decoded_lo_lo_53 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_56 , core_id_ctrl_decoder_decoded_andMatrixInput_5_56 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_55 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_20 , core_id_ctrl_decoder_decoded_andMatrixInput_6_55 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_56 , core_id_ctrl_decoder_decoded_andMatrixInput_3_56 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_39 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_56 , core_id_ctrl_decoder_decoded_andMatrixInput_1_56 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_56 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_39 , core_id_ctrl_decoder_decoded_hi_hi_lo_19 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_56 ={ core_id_ctrl_decoder_decoded_hi_hi_56 , core_id_ctrl_decoder_decoded_hi_lo_55 }; 
    wire[13:0] core__id_ctrl_decoder_decoded_T_112 ={ core_id_ctrl_decoder_decoded_hi_56 , core_id_ctrl_decoder_decoded_lo_56 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_54 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_22 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_6 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_5 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_9 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_7 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_19 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_3 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_2 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28_1 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_25 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_4 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28_2 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_6 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28_3 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_15_8 , core_id_ctrl_decoder_decoded_andMatrixInput_16_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_13_19 , core_id_ctrl_decoder_decoded_andMatrixInput_14_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_54 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_21 , core_id_ctrl_decoder_decoded_lo_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_21 , core_id_ctrl_decoder_decoded_andMatrixInput_12_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_24 , core_id_ctrl_decoder_decoded_andMatrixInput_10_21 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_57 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_24 , core_id_ctrl_decoder_decoded_lo_hi_lo_19 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_57 ={ core_id_ctrl_decoder_decoded_lo_hi_57 , core_id_ctrl_decoder_decoded_lo_lo_54 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_54 , core_id_ctrl_decoder_decoded_andMatrixInput_8_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_57 , core_id_ctrl_decoder_decoded_andMatrixInput_6_56 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_56 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_21 , core_id_ctrl_decoder_decoded_hi_lo_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_57 , core_id_ctrl_decoder_decoded_andMatrixInput_4_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_57 , core_id_ctrl_decoder_decoded_andMatrixInput_1_57 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_hi_40 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_2_57 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_hi_57 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_40 , core_id_ctrl_decoder_decoded_hi_hi_lo_20 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_hi_57 ={ core_id_ctrl_decoder_decoded_hi_hi_57 , core_id_ctrl_decoder_decoded_hi_lo_56 }; 
    wire[16:0] core__id_ctrl_decoder_decoded_T_114 ={ core_id_ctrl_decoder_decoded_hi_57 , core_id_ctrl_decoder_decoded_lo_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_2 , core_id_ctrl_decoder_decoded_andMatrixInput_19_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_15_9 , core_id_ctrl_decoder_decoded_andMatrixInput_16_3 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_hi_22 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_17_2 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_lo_55 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_22 , core_id_ctrl_decoder_decoded_lo_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_13_20 , core_id_ctrl_decoder_decoded_andMatrixInput_14_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_22 , core_id_ctrl_decoder_decoded_andMatrixInput_11_22 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_hi_25 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_12_21 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_hi_58 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_25 , core_id_ctrl_decoder_decoded_lo_hi_lo_20 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_lo_58 ={ core_id_ctrl_decoder_decoded_lo_hi_58 , core_id_ctrl_decoder_decoded_lo_lo_55 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_41 , core_id_ctrl_decoder_decoded_andMatrixInput_9_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_58 , core_id_ctrl_decoder_decoded_andMatrixInput_6_57 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_hi_22 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_7_55 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_lo_57 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_22 , core_id_ctrl_decoder_decoded_hi_lo_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_58 , core_id_ctrl_decoder_decoded_andMatrixInput_4_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_58 , core_id_ctrl_decoder_decoded_andMatrixInput_1_58 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_hi_41 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_andMatrixInput_2_58 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_hi_58 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_41 , core_id_ctrl_decoder_decoded_hi_hi_lo_21 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_hi_58 ={ core_id_ctrl_decoder_decoded_hi_hi_58 , core_id_ctrl_decoder_decoded_hi_lo_57 }; 
    wire[19:0] core__id_ctrl_decoder_decoded_T_116 ={ core_id_ctrl_decoder_decoded_hi_58 , core_id_ctrl_decoder_decoded_lo_58 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_3 = core_id_ctrl_decoder_decoded_plaInput [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_3 = core_id_ctrl_decoder_decoded_plaInput [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_3 = core_id_ctrl_decoder_decoded_plaInput [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_3 = core_id_ctrl_decoder_decoded_plaInput [22]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_25_2 , core_id_ctrl_decoder_decoded_andMatrixInput_26_2 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_10 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_27_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_23_2 , core_id_ctrl_decoder_decoded_andMatrixInput_24_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_21_2 , core_id_ctrl_decoder_decoded_andMatrixInput_22_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_23 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_56 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_23 , core_id_ctrl_decoder_decoded_lo_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_3 , core_id_ctrl_decoder_decoded_andMatrixInput_19_3 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_21 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_20_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_4 , core_id_ctrl_decoder_decoded_andMatrixInput_17_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_18 , core_id_ctrl_decoder_decoded_andMatrixInput_15_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_26 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_59 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_26 , core_id_ctrl_decoder_decoded_lo_hi_lo_21 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_59 ={ core_id_ctrl_decoder_decoded_lo_hi_59 , core_id_ctrl_decoder_decoded_lo_lo_56 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_23 , core_id_ctrl_decoder_decoded_andMatrixInput_12_22 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_18 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_13_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_26 , core_id_ctrl_decoder_decoded_andMatrixInput_10_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_56 , core_id_ctrl_decoder_decoded_andMatrixInput_8_42 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_23 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_58 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_23 , core_id_ctrl_decoder_decoded_hi_lo_lo_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_59 , core_id_ctrl_decoder_decoded_andMatrixInput_5_59 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_22 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_6_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_59 , core_id_ctrl_decoder_decoded_andMatrixInput_3_59 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_59 , core_id_ctrl_decoder_decoded_andMatrixInput_1_59 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_42 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_59 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_42 , core_id_ctrl_decoder_decoded_hi_hi_lo_22 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_59 ={ core_id_ctrl_decoder_decoded_hi_hi_59 , core_id_ctrl_decoder_decoded_hi_lo_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28_1 , core_id_ctrl_decoder_decoded_andMatrixInput_29_1 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_11 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_3 , core_id_ctrl_decoder_decoded_andMatrixInput_30_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_3 , core_id_ctrl_decoder_decoded_andMatrixInput_27_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_3 , core_id_ctrl_decoder_decoded_andMatrixInput_25_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_24 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_57 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_24 , core_id_ctrl_decoder_decoded_lo_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_3 , core_id_ctrl_decoder_decoded_andMatrixInput_23_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_3 , core_id_ctrl_decoder_decoded_andMatrixInput_21_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_22 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_4 , core_id_ctrl_decoder_decoded_andMatrixInput_19_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_5 , core_id_ctrl_decoder_decoded_andMatrixInput_17_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_27 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_60 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_27 , core_id_ctrl_decoder_decoded_lo_hi_lo_22 }; 
    wire[14:0] core_id_ctrl_decoder_decoded_lo_60 ={ core_id_ctrl_decoder_decoded_lo_hi_60 , core_id_ctrl_decoder_decoded_lo_lo_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_19 , core_id_ctrl_decoder_decoded_andMatrixInput_15_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_23 , core_id_ctrl_decoder_decoded_andMatrixInput_13_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_19 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_24 , core_id_ctrl_decoder_decoded_andMatrixInput_11_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_43 , core_id_ctrl_decoder_decoded_andMatrixInput_9_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_24 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_59 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_24 , core_id_ctrl_decoder_decoded_hi_lo_lo_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_59 , core_id_ctrl_decoder_decoded_andMatrixInput_7_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_60 , core_id_ctrl_decoder_decoded_andMatrixInput_5_60 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_23 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_60 , core_id_ctrl_decoder_decoded_andMatrixInput_3_60 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_60 , core_id_ctrl_decoder_decoded_andMatrixInput_1_60 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_43 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_60 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_43 , core_id_ctrl_decoder_decoded_hi_hi_lo_23 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_60 ={ core_id_ctrl_decoder_decoded_hi_hi_60 , core_id_ctrl_decoder_decoded_hi_lo_59 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_24 , core_id_ctrl_decoder_decoded_andMatrixInput_13_23 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_58 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_25 , core_id_ctrl_decoder_decoded_andMatrixInput_14_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_25 , core_id_ctrl_decoder_decoded_andMatrixInput_11_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_44 , core_id_ctrl_decoder_decoded_andMatrixInput_9_28 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_61 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_28 , core_id_ctrl_decoder_decoded_lo_hi_lo_23 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_61 ={ core_id_ctrl_decoder_decoded_lo_hi_61 , core_id_ctrl_decoder_decoded_lo_lo_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_60 , core_id_ctrl_decoder_decoded_andMatrixInput_7_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_61 , core_id_ctrl_decoder_decoded_andMatrixInput_5_61 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_60 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_25 , core_id_ctrl_decoder_decoded_hi_lo_lo_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_61 , core_id_ctrl_decoder_decoded_andMatrixInput_3_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_61 , core_id_ctrl_decoder_decoded_andMatrixInput_1_61 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_61 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_44 , core_id_ctrl_decoder_decoded_hi_hi_lo_24 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_61 ={ core_id_ctrl_decoder_decoded_hi_hi_61 , core_id_ctrl_decoder_decoded_hi_lo_60 }; 
    wire[14:0] core__id_ctrl_decoder_decoded_T_122 ={ core_id_ctrl_decoder_decoded_hi_61 , core_id_ctrl_decoder_decoded_lo_61 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_25 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_4 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29_2 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_6 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29_3 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_26 , core_id_ctrl_decoder_decoded_andMatrixInput_11_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_59 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_26 , core_id_ctrl_decoder_decoded_andMatrixInput_12_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_59 , core_id_ctrl_decoder_decoded_andMatrixInput_8_45 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_62 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_29 , core_id_ctrl_decoder_decoded_andMatrixInput_9_29 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_62 ={ core_id_ctrl_decoder_decoded_lo_hi_62 , core_id_ctrl_decoder_decoded_lo_lo_59 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_62 , core_id_ctrl_decoder_decoded_andMatrixInput_5_62 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_61 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_26 , core_id_ctrl_decoder_decoded_andMatrixInput_6_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_62 , core_id_ctrl_decoder_decoded_andMatrixInput_3_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_45 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_62 , core_id_ctrl_decoder_decoded_andMatrixInput_1_62 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_62 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_45 , core_id_ctrl_decoder_decoded_hi_hi_lo_25 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_62 ={ core_id_ctrl_decoder_decoded_hi_hi_62 , core_id_ctrl_decoder_decoded_hi_lo_61 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_5 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_5 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_7 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_7 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_25_4 , core_id_ctrl_decoder_decoded_andMatrixInput_26_4 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_12 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_27_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_23_4 , core_id_ctrl_decoder_decoded_andMatrixInput_24_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_21_4 , core_id_ctrl_decoder_decoded_andMatrixInput_22_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_27 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_60 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_27 , core_id_ctrl_decoder_decoded_lo_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_5 , core_id_ctrl_decoder_decoded_andMatrixInput_19_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_24 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_20_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_6 , core_id_ctrl_decoder_decoded_andMatrixInput_17_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_21 , core_id_ctrl_decoder_decoded_andMatrixInput_15_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_30 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_63 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_30 , core_id_ctrl_decoder_decoded_lo_hi_lo_24 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_63 ={ core_id_ctrl_decoder_decoded_lo_hi_63 , core_id_ctrl_decoder_decoded_lo_lo_60 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_27 , core_id_ctrl_decoder_decoded_andMatrixInput_12_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_21 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_13_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_30 , core_id_ctrl_decoder_decoded_andMatrixInput_10_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_60 , core_id_ctrl_decoder_decoded_andMatrixInput_8_46 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_27 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_62 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_27 , core_id_ctrl_decoder_decoded_hi_lo_lo_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_63 , core_id_ctrl_decoder_decoded_andMatrixInput_5_63 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_26 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_6_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_63 , core_id_ctrl_decoder_decoded_andMatrixInput_3_63 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_63 , core_id_ctrl_decoder_decoded_andMatrixInput_1_63 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_46 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_63 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_46 , core_id_ctrl_decoder_decoded_hi_hi_lo_26 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_63 ={ core_id_ctrl_decoder_decoded_hi_hi_63 , core_id_ctrl_decoder_decoded_hi_lo_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_30_2 , core_id_ctrl_decoder_decoded_andMatrixInput_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28_2 , core_id_ctrl_decoder_decoded_andMatrixInput_29_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_lo_13 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_5 , core_id_ctrl_decoder_decoded_andMatrixInput_27_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_5 , core_id_ctrl_decoder_decoded_andMatrixInput_25_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_28 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_lo_61 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_28 , core_id_ctrl_decoder_decoded_lo_lo_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_5 , core_id_ctrl_decoder_decoded_andMatrixInput_23_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_5 , core_id_ctrl_decoder_decoded_andMatrixInput_21_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_25 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_6 , core_id_ctrl_decoder_decoded_andMatrixInput_19_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_7 , core_id_ctrl_decoder_decoded_andMatrixInput_17_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_31 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_64 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_31 , core_id_ctrl_decoder_decoded_lo_hi_lo_25 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_lo_64 ={ core_id_ctrl_decoder_decoded_lo_hi_64 , core_id_ctrl_decoder_decoded_lo_lo_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_22 , core_id_ctrl_decoder_decoded_andMatrixInput_15_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_27 , core_id_ctrl_decoder_decoded_andMatrixInput_13_25 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_22 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_28 , core_id_ctrl_decoder_decoded_andMatrixInput_11_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_47 , core_id_ctrl_decoder_decoded_andMatrixInput_9_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_28 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_63 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_28 , core_id_ctrl_decoder_decoded_hi_lo_lo_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_63 , core_id_ctrl_decoder_decoded_andMatrixInput_7_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_64 , core_id_ctrl_decoder_decoded_andMatrixInput_5_64 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_27 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_64 , core_id_ctrl_decoder_decoded_andMatrixInput_3_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_64 , core_id_ctrl_decoder_decoded_andMatrixInput_1_64 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_47 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_64 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_47 , core_id_ctrl_decoder_decoded_hi_hi_lo_27 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_64 ={ core_id_ctrl_decoder_decoded_hi_hi_64 , core_id_ctrl_decoder_decoded_hi_lo_63 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_14 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_29 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_24 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_6 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30_3 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_15_14 , core_id_ctrl_decoder_decoded_andMatrixInput_16_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_13_26 , core_id_ctrl_decoder_decoded_andMatrixInput_14_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_62 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_29 , core_id_ctrl_decoder_decoded_lo_lo_lo_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_29 , core_id_ctrl_decoder_decoded_andMatrixInput_12_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_32 , core_id_ctrl_decoder_decoded_andMatrixInput_10_29 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_65 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_32 , core_id_ctrl_decoder_decoded_lo_hi_lo_26 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_65 ={ core_id_ctrl_decoder_decoded_lo_hi_65 , core_id_ctrl_decoder_decoded_lo_lo_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_62 , core_id_ctrl_decoder_decoded_andMatrixInput_8_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_65 , core_id_ctrl_decoder_decoded_andMatrixInput_6_64 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_64 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_29 , core_id_ctrl_decoder_decoded_hi_lo_lo_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_65 , core_id_ctrl_decoder_decoded_andMatrixInput_4_65 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_65 , core_id_ctrl_decoder_decoded_andMatrixInput_1_65 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_hi_48 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_andMatrixInput_2_65 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_hi_65 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_48 , core_id_ctrl_decoder_decoded_hi_hi_lo_28 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_hi_65 ={ core_id_ctrl_decoder_decoded_hi_hi_65 , core_id_ctrl_decoder_decoded_hi_lo_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_30 , core_id_ctrl_decoder_decoded_andMatrixInput_11_30 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_63 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_30 , core_id_ctrl_decoder_decoded_andMatrixInput_12_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_63 , core_id_ctrl_decoder_decoded_andMatrixInput_8_49 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_66 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_33 , core_id_ctrl_decoder_decoded_andMatrixInput_9_33 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_66 ={ core_id_ctrl_decoder_decoded_lo_hi_66 , core_id_ctrl_decoder_decoded_lo_lo_63 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_66 , core_id_ctrl_decoder_decoded_andMatrixInput_5_66 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_65 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_30 , core_id_ctrl_decoder_decoded_andMatrixInput_6_65 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_66 , core_id_ctrl_decoder_decoded_andMatrixInput_3_66 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_66 , core_id_ctrl_decoder_decoded_andMatrixInput_1_66 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_66 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_49 , core_id_ctrl_decoder_decoded_hi_hi_lo_29 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_66 ={ core_id_ctrl_decoder_decoded_hi_hi_66 , core_id_ctrl_decoder_decoded_hi_lo_65 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_24 , core_id_ctrl_decoder_decoded_andMatrixInput_15_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_30 , core_id_ctrl_decoder_decoded_andMatrixInput_13_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_64 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_31 , core_id_ctrl_decoder_decoded_lo_lo_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_31 , core_id_ctrl_decoder_decoded_andMatrixInput_11_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_50 , core_id_ctrl_decoder_decoded_andMatrixInput_9_34 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_67 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_34 , core_id_ctrl_decoder_decoded_lo_hi_lo_27 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_67 ={ core_id_ctrl_decoder_decoded_lo_hi_67 , core_id_ctrl_decoder_decoded_lo_lo_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_66 , core_id_ctrl_decoder_decoded_andMatrixInput_7_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_67 , core_id_ctrl_decoder_decoded_andMatrixInput_5_67 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_66 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_31 , core_id_ctrl_decoder_decoded_hi_lo_lo_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_67 , core_id_ctrl_decoder_decoded_andMatrixInput_3_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_50 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_67 , core_id_ctrl_decoder_decoded_andMatrixInput_1_67 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_67 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_50 , core_id_ctrl_decoder_decoded_hi_hi_lo_30 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_67 ={ core_id_ctrl_decoder_decoded_hi_hi_67 , core_id_ctrl_decoder_decoded_hi_lo_66 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_6 = core_id_ctrl_decoder_decoded_plaInput [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_7 = core_id_ctrl_decoder_decoded_plaInput [24]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_25_6 , core_id_ctrl_decoder_decoded_andMatrixInput_26_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_16 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_27_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_23_6 , core_id_ctrl_decoder_decoded_andMatrixInput_24_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_21_6 , core_id_ctrl_decoder_decoded_andMatrixInput_22_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_32 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_65 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_32 , core_id_ctrl_decoder_decoded_lo_lo_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_7 , core_id_ctrl_decoder_decoded_andMatrixInput_19_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_28 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_20_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_9 , core_id_ctrl_decoder_decoded_andMatrixInput_17_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_25 , core_id_ctrl_decoder_decoded_andMatrixInput_15_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_35 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_68 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_35 , core_id_ctrl_decoder_decoded_lo_hi_lo_28 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_68 ={ core_id_ctrl_decoder_decoded_lo_hi_68 , core_id_ctrl_decoder_decoded_lo_lo_65 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_32 , core_id_ctrl_decoder_decoded_andMatrixInput_12_31 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_25 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_13_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_35 , core_id_ctrl_decoder_decoded_andMatrixInput_10_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_65 , core_id_ctrl_decoder_decoded_andMatrixInput_8_51 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_32 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_67 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_32 , core_id_ctrl_decoder_decoded_hi_lo_lo_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_68 , core_id_ctrl_decoder_decoded_andMatrixInput_5_68 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_31 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_6_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_68 , core_id_ctrl_decoder_decoded_andMatrixInput_3_68 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_68 , core_id_ctrl_decoder_decoded_andMatrixInput_1_68 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_51 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_9 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_68 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_51 , core_id_ctrl_decoder_decoded_hi_hi_lo_31 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_68 ={ core_id_ctrl_decoder_decoded_hi_hi_68 , core_id_ctrl_decoder_decoded_hi_lo_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_30_3 , core_id_ctrl_decoder_decoded_andMatrixInput_31_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28_3 , core_id_ctrl_decoder_decoded_andMatrixInput_29_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_lo_17 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_lo_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_7 , core_id_ctrl_decoder_decoded_andMatrixInput_27_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_7 , core_id_ctrl_decoder_decoded_andMatrixInput_25_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_33 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_8 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_lo_66 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_33 , core_id_ctrl_decoder_decoded_lo_lo_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_7 , core_id_ctrl_decoder_decoded_andMatrixInput_23_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_7 , core_id_ctrl_decoder_decoded_andMatrixInput_21_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_29 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_8 , core_id_ctrl_decoder_decoded_andMatrixInput_19_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_10 , core_id_ctrl_decoder_decoded_andMatrixInput_17_8 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_36 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_69 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_36 , core_id_ctrl_decoder_decoded_lo_hi_lo_29 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_lo_69 ={ core_id_ctrl_decoder_decoded_lo_hi_69 , core_id_ctrl_decoder_decoded_lo_lo_66 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_26 , core_id_ctrl_decoder_decoded_andMatrixInput_15_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_32 , core_id_ctrl_decoder_decoded_andMatrixInput_13_29 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_26 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_33 , core_id_ctrl_decoder_decoded_andMatrixInput_11_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_52 , core_id_ctrl_decoder_decoded_andMatrixInput_9_36 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_33 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_8 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_68 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_33 , core_id_ctrl_decoder_decoded_hi_lo_lo_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_68 , core_id_ctrl_decoder_decoded_andMatrixInput_7_66 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_69 , core_id_ctrl_decoder_decoded_andMatrixInput_5_69 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_32 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_69 , core_id_ctrl_decoder_decoded_andMatrixInput_3_69 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_69 , core_id_ctrl_decoder_decoded_andMatrixInput_1_69 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_52 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_10 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_69 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_52 , core_id_ctrl_decoder_decoded_hi_hi_lo_32 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_69 ={ core_id_ctrl_decoder_decoded_hi_hi_69 , core_id_ctrl_decoder_decoded_hi_lo_68 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_33 = core_id_ctrl_decoder_decoded_plaInput [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_34 , core_id_ctrl_decoder_decoded_andMatrixInput_11_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_67 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_34 , core_id_ctrl_decoder_decoded_andMatrixInput_12_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_67 , core_id_ctrl_decoder_decoded_andMatrixInput_8_53 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_70 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_37 , core_id_ctrl_decoder_decoded_andMatrixInput_9_37 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_70 ={ core_id_ctrl_decoder_decoded_lo_hi_70 , core_id_ctrl_decoder_decoded_lo_lo_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_70 , core_id_ctrl_decoder_decoded_andMatrixInput_5_70 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_69 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_34 , core_id_ctrl_decoder_decoded_andMatrixInput_6_69 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_70 , core_id_ctrl_decoder_decoded_andMatrixInput_3_70 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_53 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_70 , core_id_ctrl_decoder_decoded_andMatrixInput_1_70 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_70 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_53 , core_id_ctrl_decoder_decoded_hi_hi_lo_33 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_70 ={ core_id_ctrl_decoder_decoded_hi_hi_70 , core_id_ctrl_decoder_decoded_hi_lo_69 }; 
    wire[1:0] core__GEN_0 ={& core__id_ctrl_decoder_decoded_T_58 ,& core__id_ctrl_decoder_decoded_T_112 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi = core__GEN_0 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_2 = core__GEN_0 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi ={&{ core_id_ctrl_decoder_decoded_hi_59 , core_id_ctrl_decoder_decoded_lo_59 },&{ core_id_ctrl_decoder_decoded_hi_63 , core_id_ctrl_decoder_decoded_lo_63 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi ,&{ core_id_ctrl_decoder_decoded_hi_68 , core_id_ctrl_decoder_decoded_lo_68 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi ={&{ core_id_ctrl_decoder_decoded_hi_18 , core_id_ctrl_decoder_decoded_lo_18 },& core__id_ctrl_decoder_decoded_T_52 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi ,& core__id_ctrl_decoder_decoded_T_64 }; 
    wire[1:0] core__GEN_1 ={& core__id_ctrl_decoder_decoded_T_112 ,& core__id_ctrl_decoder_decoded_T_114 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo = core__GEN_1 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_5 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_5 = core__GEN_1 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_1 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_1 = core__GEN_1 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_2 = core__GEN_1 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_3 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_3 = core__GEN_1 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_8 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_8 = core__GEN_1 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi ={& core__id_ctrl_decoder_decoded_T_64 ,& core__id_ctrl_decoder_decoded_T_78 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo ={& core__id_ctrl_decoder_decoded_T_54 ,& core__id_ctrl_decoder_decoded_T_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi ={& core__id_ctrl_decoder_decoded_T_42 ,& core__id_ctrl_decoder_decoded_T_52 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo }; 
    wire[7:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo ={& core__id_ctrl_decoder_decoded_T_32 ,& core__id_ctrl_decoder_decoded_T_34 }; 
    wire[1:0] core__GEN_2 ={& core__id_ctrl_decoder_decoded_T_22 ,& core__id_ctrl_decoder_decoded_T_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi = core__GEN_2 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_1 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_1 = core__GEN_2 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_2 = core__GEN_2 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_5 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_5 = core__GEN_2 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi = core__GEN_2 ; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo ={& core__id_ctrl_decoder_decoded_T_6 ,& core__id_ctrl_decoder_decoded_T_12 }; 
    wire[1:0] core__GEN_3 ={& core__id_ctrl_decoder_decoded_T ,&{ core_id_ctrl_decoder_decoded_hi_1 , core_id_ctrl_decoder_decoded_lo_1 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_3 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_3 = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_4 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_4 = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_5 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_5 = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_6 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_6 = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_7 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_7 = core__GEN_3 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_1 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_1 = core__GEN_3 ; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo }; 
    wire[7:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_2 ={& core__id_ctrl_decoder_decoded_T_122 ,&{ core_id_ctrl_decoder_decoded_hi_62 , core_id_ctrl_decoder_decoded_lo_62 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_3 ={& core__id_ctrl_decoder_decoded_T_16 ,&{ core_id_ctrl_decoder_decoded_hi_10 , core_id_ctrl_decoder_decoded_lo_10 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_4 ={& core__id_ctrl_decoder_decoded_T_114 ,& core__id_ctrl_decoder_decoded_T_122 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_2 ,& core__id_ctrl_decoder_decoded_T_116 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_2 ={& core__id_ctrl_decoder_decoded_T ,& core__id_ctrl_decoder_decoded_T_4 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_2 ,& core__id_ctrl_decoder_decoded_T_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_3 ={&{ core_id_ctrl_decoder_decoded_hi_45 , core_id_ctrl_decoder_decoded_lo_45 },&{ core_id_ctrl_decoder_decoded_hi_52 , core_id_ctrl_decoder_decoded_lo_52 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_3 ,&{ core_id_ctrl_decoder_decoded_hi_54 , core_id_ctrl_decoder_decoded_lo_54 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_1 ={& core__id_ctrl_decoder_decoded_T_78 ,&{ core_id_ctrl_decoder_decoded_hi_43 , core_id_ctrl_decoder_decoded_lo_43 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_3 ={& core__id_ctrl_decoder_decoded_T_42 ,&{ core_id_ctrl_decoder_decoded_hi_24 , core_id_ctrl_decoder_decoded_lo_24 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_1 }; 
    wire[1:0] core__GEN_4 ={&{ core_id_ctrl_decoder_decoded_hi_65 , core_id_ctrl_decoder_decoded_lo_65 },&{ core_id_ctrl_decoder_decoded_hi_67 , core_id_ctrl_decoder_decoded_lo_67 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_1 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_1 = core__GEN_4 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_7 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_7 = core__GEN_4 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_4 ={&{ core_id_ctrl_decoder_decoded_hi_50 , core_id_ctrl_decoder_decoded_lo_50 },&{ core_id_ctrl_decoder_decoded_hi_55 , core_id_ctrl_decoder_decoded_lo_55 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_2 ={&{ core_id_ctrl_decoder_decoded_hi_47 , core_id_ctrl_decoder_decoded_lo_47 },&{ core_id_ctrl_decoder_decoded_hi_48 , core_id_ctrl_decoder_decoded_lo_48 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_1 ={&{ core_id_ctrl_decoder_decoded_hi_14 , core_id_ctrl_decoder_decoded_lo_14 },&{ core_id_ctrl_decoder_decoded_hi_34 , core_id_ctrl_decoder_decoded_lo_34 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_1 ,&{ core_id_ctrl_decoder_decoded_hi_35 , core_id_ctrl_decoder_decoded_lo_35 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_5 ={&{ core_id_ctrl_decoder_decoded_hi_37 , core_id_ctrl_decoder_decoded_lo_37 },& core__id_ctrl_decoder_decoded_T_76 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_5 ,&{ core_id_ctrl_decoder_decoded_hi_41 , core_id_ctrl_decoder_decoded_lo_41 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_5 ={& core__id_ctrl_decoder_decoded_T_54 ,&{ core_id_ctrl_decoder_decoded_hi_30 , core_id_ctrl_decoder_decoded_lo_30 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_5 ,&{ core_id_ctrl_decoder_decoded_hi_36 , core_id_ctrl_decoder_decoded_lo_36 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_6 ={&{ core_id_ctrl_decoder_decoded_hi_28 , core_id_ctrl_decoder_decoded_lo_28 },&{ core_id_ctrl_decoder_decoded_hi_31 , core_id_ctrl_decoder_decoded_lo_31 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_6 ,& core__id_ctrl_decoder_decoded_T_76 }; 
    wire[1:0] core__GEN_5 ={& core__id_ctrl_decoder_decoded_T_76 ,& core__id_ctrl_decoder_decoded_T_78 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_1 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_1 = core__GEN_5 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_2 = core__GEN_5 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_5 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_5 = core__GEN_5 ; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_1 ={& core__id_ctrl_decoder_decoded_T_58 ,& core__id_ctrl_decoder_decoded_T_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi ={& core__id_ctrl_decoder_decoded_T_42 ,& core__id_ctrl_decoder_decoded_T_46 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi ,& core__id_ctrl_decoder_decoded_T_54 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_1 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_1 ={& core__id_ctrl_decoder_decoded_T_30 ,& core__id_ctrl_decoder_decoded_T_34 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_1 }; 
    wire[1:0] core__GEN_6 ={& core__id_ctrl_decoder_decoded_T_8 ,& core__id_ctrl_decoder_decoded_T_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_1 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_1 = core__GEN_6 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_3 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_3 = core__GEN_6 ; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi ,& core__id_ctrl_decoder_decoded_T_4 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_1 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_9 ={& core__id_ctrl_decoder_decoded_T_88 ,& core__id_ctrl_decoder_decoded_T_98 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_12 ={& core__id_ctrl_decoder_decoded_T_26 ,& core__id_ctrl_decoder_decoded_T_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_3 ={& core__id_ctrl_decoder_decoded_T_92 ,& core__id_ctrl_decoder_decoded_T_102 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_7 ={& core__id_ctrl_decoder_decoded_T_54 ,& core__id_ctrl_decoder_decoded_T_80 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_4 ={& core__id_ctrl_decoder_decoded_T_32 ,& core__id_ctrl_decoder_decoded_T_44 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_3 ,& core__id_ctrl_decoder_decoded_T_6 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_2 }; 
    wire[1:0] core__GEN_7 ={& core__id_ctrl_decoder_decoded_T_58 ,&{ core_id_ctrl_decoder_decoded_hi_33 , core_id_ctrl_decoder_decoded_lo_33 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_2 = core__GEN_7 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_4 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_4 = core__GEN_7 ; 
    wire[1:0] core__GEN_8 ={&{ core_id_ctrl_decoder_decoded_hi_25 , core_id_ctrl_decoder_decoded_lo_25 },& core__id_ctrl_decoder_decoded_T_54 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_2 = core__GEN_8 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_5 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_5 = core__GEN_8 ; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_2 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_4 }; 
    wire[1:0] core__GEN_9 ={& core__id_ctrl_decoder_decoded_T_30 ,& core__id_ctrl_decoder_decoded_T_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_2 = core__GEN_9 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_3 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_3 = core__GEN_9 ; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_2 }; 
    wire[1:0] core__GEN_10 ={& core__id_ctrl_decoder_decoded_T_4 ,& core__id_ctrl_decoder_decoded_T_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_2 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_2 = core__GEN_10 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_3 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_3 = core__GEN_10 ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_4 ; 
  assign  core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_4 = core__GEN_10 ; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_2 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_3 ={& core__id_ctrl_decoder_decoded_T_80 ,& core__id_ctrl_decoder_decoded_T_92 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_3 ,& core__id_ctrl_decoder_decoded_T_102 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_3 ={& core__id_ctrl_decoder_decoded_T_34 ,& core__id_ctrl_decoder_decoded_T_44 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_3 ,& core__id_ctrl_decoder_decoded_T_54 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_3 ,& core__id_ctrl_decoder_decoded_T_32 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_5 ,& core__id_ctrl_decoder_decoded_T_4 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_4 ={& core__id_ctrl_decoder_decoded_T_78 ,& core__id_ctrl_decoder_decoded_T_88 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_4 ,& core__id_ctrl_decoder_decoded_T_98 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_3 ={& core__id_ctrl_decoder_decoded_T_42 ,& core__id_ctrl_decoder_decoded_T_54 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_4 ={& core__id_ctrl_decoder_decoded_T_26 ,& core__id_ctrl_decoder_decoded_T_30 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_4 ={& core__id_ctrl_decoder_decoded_T_12 ,& core__id_ctrl_decoder_decoded_T_22 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_4 ,& core__id_ctrl_decoder_decoded_T_24 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_16 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_4 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_4 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_17 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_12 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_12 ={& core__id_ctrl_decoder_decoded_T_76 ,&{ core_id_ctrl_decoder_decoded_hi_42 , core_id_ctrl_decoder_decoded_lo_42 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_12 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_9 ={& core__id_ctrl_decoder_decoded_T_24 ,& core__id_ctrl_decoder_decoded_T_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_8 ={& core__id_ctrl_decoder_decoded_T_16 ,&{ core_id_ctrl_decoder_decoded_hi_9 , core_id_ctrl_decoder_decoded_lo_9 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_8 ,& core__id_ctrl_decoder_decoded_T_22 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_18 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_13 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_4 ={&{ core_id_ctrl_decoder_decoded_hi_64 , core_id_ctrl_decoder_decoded_lo_64 },&{ core_id_ctrl_decoder_decoded_hi_69 , core_id_ctrl_decoder_decoded_lo_69 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi ={& core__id_ctrl_decoder_decoded_T_112 ,& core__id_ctrl_decoder_decoded_T_116 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi ,&{ core_id_ctrl_decoder_decoded_hi_60 , core_id_ctrl_decoder_decoded_lo_60 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi ={& core__id_ctrl_decoder_decoded_T_64 ,& core__id_ctrl_decoder_decoded_T_76 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi ,& core__id_ctrl_decoder_decoded_T_78 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_1 ={& core__id_ctrl_decoder_decoded_T_46 ,& core__id_ctrl_decoder_decoded_T_54 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_1 ,& core__id_ctrl_decoder_decoded_T_58 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_5 }; 
    wire[10:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_16 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_13 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi ={& core__id_ctrl_decoder_decoded_T_34 ,&{ core_id_ctrl_decoder_decoded_hi_19 , core_id_ctrl_decoder_decoded_lo_19 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi ,& core__id_ctrl_decoder_decoded_T_42 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi ,& core__id_ctrl_decoder_decoded_T_30 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi ={& core__id_ctrl_decoder_decoded_T_8 ,& core__id_ctrl_decoder_decoded_T_10 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi ,& core__id_ctrl_decoder_decoded_T_12 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_1 ,& core__id_ctrl_decoder_decoded_T_4 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_5 }; 
    wire[11:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_19 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_14 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi ,& core__id_ctrl_decoder_decoded_T_114 },1'h0}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi_hi ={& core__id_ctrl_decoder_decoded_T_52 ,&{ core_id_ctrl_decoder_decoded_hi_20 , core_id_ctrl_decoder_decoded_lo_20 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi_hi ,& core__id_ctrl_decoder_decoded_T_10 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo },& core__id_ctrl_decoder_decoded_T_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_hi ={1'h0,&{ core_id_ctrl_decoder_decoded_hi_53 , core_id_ctrl_decoder_decoded_lo_53 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_1 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_2 },1'h0}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_hi ,1'h0}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_1 ,2'h0}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_5 ,&{ core_id_ctrl_decoder_decoded_hi_70 , core_id_ctrl_decoder_decoded_lo_70 }},|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_4 ,&{ core_id_ctrl_decoder_decoded_hi_66 , core_id_ctrl_decoder_decoded_lo_66 }}}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_3 },1'h0}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_hi ,& core__id_ctrl_decoder_decoded_T_58 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_6 }; 
    wire[19:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_17 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_14 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_5 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_4 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_8 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_7 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_6 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_lo ={|{& core__id_ctrl_decoder_decoded_T_12 ,& core__id_ctrl_decoder_decoded_T_34 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_12 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_9 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_hi ={|{&{ core_id_ctrl_decoder_decoded_hi_7 , core_id_ctrl_decoder_decoded_lo_7 },& core__id_ctrl_decoder_decoded_T_34 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_14 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_11 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_13 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_10 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_16 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_13 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_15 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_12 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_hi ={& core__id_ctrl_decoder_decoded_T_32 ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_18 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_15 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_17 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_14 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_lo ={|{& core__id_ctrl_decoder_decoded_T_26 ,& core__id_ctrl_decoder_decoded_T_76 },& core__id_ctrl_decoder_decoded_T_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_19 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_16 },1'h0}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_hi ,1'h0}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6 }; 
    wire[19:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_20 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_15 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_11 }; 
    wire[39:0] core_id_ctrl_decoder_decoded_orMatrixOutputs ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_20 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [1:0]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [4:3]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [2]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [6:5]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [9:8]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [7]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [11:10]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [14:13]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [12]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [16:15]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [19:18]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [17]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo }; 
    wire[19:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [21:20]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [24:23]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [22]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [26:25]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [29:28]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [27]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [31:30]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [34:33]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [32]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_lo = core_id_ctrl_decoder_decoded_orMatrixOutputs [36:35]; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi_hi = core_id_ctrl_decoder_decoded_orMatrixOutputs [39:38]; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [37]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo }; 
    wire[19:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo }; 
  assign  core_id_ctrl_decoder_decoded_invMatrixOutputs ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo }; 
    wire[39:0] core_id_ctrl_decoder_decoded = core_id_ctrl_decoder_decoded_invMatrixOutputs ; 
  assign  core_id_ctrl_decoder_0 = core_id_ctrl_decoder_decoded [39]; 
    wire core_id_ctrl_legal = core_id_ctrl_decoder_0 ; 
  assign  core_id_ctrl_decoder_1 = core_id_ctrl_decoder_decoded [38]; 
    wire core_id_ctrl_fp = core_id_ctrl_decoder_1 ; 
  assign  core_id_ctrl_decoder_2 = core_id_ctrl_decoder_decoded [37]; 
    wire core_id_ctrl_rocc = core_id_ctrl_decoder_2 ; 
  assign  core_id_ctrl_decoder_3 = core_id_ctrl_decoder_decoded [36]; 
    wire core_id_ctrl_branch = core_id_ctrl_decoder_3 ; 
  assign  core_id_ctrl_decoder_4 = core_id_ctrl_decoder_decoded [35]; 
    wire core_id_ctrl_jal = core_id_ctrl_decoder_4 ; 
  assign  core_id_ctrl_decoder_5 = core_id_ctrl_decoder_decoded [34]; 
    wire core_id_ctrl_jalr = core_id_ctrl_decoder_5 ; 
  assign  core_id_ctrl_decoder_6 = core_id_ctrl_decoder_decoded [33]; 
    wire core_id_ctrl_rxs2 = core_id_ctrl_decoder_6 ; 
  assign  core_id_ctrl_decoder_7 = core_id_ctrl_decoder_decoded [32]; 
    wire core_id_ctrl_rxs1 = core_id_ctrl_decoder_7 ; 
  assign  core_id_ctrl_decoder_8 = core_id_ctrl_decoder_decoded [31:30]; 
    wire[1:0] core_id_ctrl_sel_alu2 = core_id_ctrl_decoder_8 ; 
  assign  core_id_ctrl_decoder_9 = core_id_ctrl_decoder_decoded [29:28]; 
    wire[1:0] core_id_ctrl_sel_alu1 = core_id_ctrl_decoder_9 ; 
  assign  core_id_ctrl_decoder_10 = core_id_ctrl_decoder_decoded [27:25]; 
    wire[2:0] core_id_ctrl_sel_imm = core_id_ctrl_decoder_10 ; 
  assign  core_id_ctrl_decoder_11 = core_id_ctrl_decoder_decoded [24]; 
    wire core_id_ctrl_alu_dw = core_id_ctrl_decoder_11 ; 
  assign  core_id_ctrl_decoder_12 = core_id_ctrl_decoder_decoded [23:20]; 
    wire[3:0] core_id_ctrl_alu_fn = core_id_ctrl_decoder_12 ; 
  assign  core_id_ctrl_decoder_13 = core_id_ctrl_decoder_decoded [19]; 
    wire core_id_ctrl_mem = core_id_ctrl_decoder_13 ; 
  assign  core_id_ctrl_decoder_14 = core_id_ctrl_decoder_decoded [18:14]; 
    wire[4:0] core_id_ctrl_mem_cmd = core_id_ctrl_decoder_14 ; 
  assign  core_id_ctrl_decoder_15 = core_id_ctrl_decoder_decoded [13]; 
    wire core_id_ctrl_rfs1 = core_id_ctrl_decoder_15 ; 
  assign  core_id_ctrl_decoder_16 = core_id_ctrl_decoder_decoded [12]; 
    wire core_id_ctrl_rfs2 = core_id_ctrl_decoder_16 ; 
  assign  core_id_ctrl_decoder_17 = core_id_ctrl_decoder_decoded [11]; 
    wire core_id_ctrl_rfs3 = core_id_ctrl_decoder_17 ; 
  assign  core_id_ctrl_decoder_18 = core_id_ctrl_decoder_decoded [10]; 
    wire core_id_ctrl_wfd = core_id_ctrl_decoder_18 ; 
  assign  core_id_ctrl_decoder_19 = core_id_ctrl_decoder_decoded [9]; 
    wire core_id_ctrl_mul = core_id_ctrl_decoder_19 ; 
  assign  core_id_ctrl_decoder_20 = core_id_ctrl_decoder_decoded [8]; 
    wire core_id_ctrl_div = core_id_ctrl_decoder_20 ; 
  assign  core_id_ctrl_decoder_21 = core_id_ctrl_decoder_decoded [7]; 
    wire core_id_ctrl_wxd = core_id_ctrl_decoder_21 ; 
  assign  core_id_ctrl_decoder_22 = core_id_ctrl_decoder_decoded [6:4]; 
    wire[2:0] core_id_ctrl_csr = core_id_ctrl_decoder_22 ; 
  assign  core_id_ctrl_decoder_23 = core_id_ctrl_decoder_decoded [3]; 
    wire core_id_ctrl_fence_i = core_id_ctrl_decoder_23 ; 
  assign  core_id_ctrl_decoder_24 = core_id_ctrl_decoder_decoded [2]; 
    wire core_id_ctrl_fence = core_id_ctrl_decoder_24 ; 
  assign  core_id_ctrl_decoder_25 = core_id_ctrl_decoder_decoded [1]; 
    wire core_id_ctrl_amo = core_id_ctrl_decoder_25 ; 
  assign  core_id_ctrl_decoder_26 = core_id_ctrl_decoder_decoded [0]; 
    wire core_id_ctrl_dp = core_id_ctrl_decoder_26 ; 
    reg core_id_reg_fence ; 
    wire[4:0] core_id_raddr1 ; 
    wire[4:0] core_id_raddr2 ; 
    wire core_id_npc_sign = core__ibuf_io_inst_0_bits_inst_bits [31]; 
    wire core_id_npc_hi_hi_hi = core_id_npc_sign ; 
    wire[10:0] core_id_npc_b30_20 ={11{ core_id_npc_sign }}; 
    wire[10:0] core_id_npc_hi_hi_lo = core_id_npc_b30_20 ; 
    wire[7:0] core_id_npc_b19_12 = core__ibuf_io_inst_0_bits_inst_bits [19:12]; 
    wire[7:0] core_id_npc_hi_lo_hi = core_id_npc_b19_12 ; 
    wire core_id_npc_b11 = core__ibuf_io_inst_0_bits_inst_bits [20]; 
    wire core_id_npc_hi_lo_lo = core_id_npc_b11 ; 
    wire[5:0] core_id_npc_b10_5 = core__ibuf_io_inst_0_bits_inst_bits [30:25]; 
    wire[3:0] core_id_npc_b4_1 = core__ibuf_io_inst_0_bits_inst_bits [24:21]; 
    wire[9:0] core_id_npc_lo_hi ={ core_id_npc_b10_5 , core_id_npc_b4_1 }; 
    wire[10:0] core_id_npc_lo ={ core_id_npc_lo_hi ,1'h0}; 
    wire[8:0] core_id_npc_hi_lo ={ core_id_npc_hi_lo_hi , core_id_npc_hi_lo_lo }; 
    wire[11:0] core_id_npc_hi_hi ={ core_id_npc_hi_hi_hi , core_id_npc_hi_hi_lo }; 
    wire[20:0] core_id_npc_hi ={ core_id_npc_hi_hi , core_id_npc_hi_lo }; 
    wire[31:0] core_id_npc = core__ibuf_io_pc +{ core_id_npc_hi , core_id_npc_lo }; 
    wire core__id_csr_ren_T = core_id_ctrl_csr ==3'h6; 
    wire core_id_csr_en = core__id_csr_ren_T |(& core_id_ctrl_csr )| core_id_ctrl_csr ==3'h5; 
    wire core_id_system_insn = core_id_ctrl_csr ==3'h4; 
    wire core_id_csr_ren =( core__id_csr_ren_T |(& core_id_ctrl_csr ))& core__ibuf_io_inst_0_bits_inst_rs1 ==5'h0; 
    wire[2:0] core_id_csr = core_id_system_insn & core_id_ctrl_mem  ? 3'h0: core_id_csr_ren  ? 3'h2: core_id_ctrl_csr ; 
    wire core_id_csr_flush = core_id_system_insn | core_id_csr_en &~ core_id_csr_ren & core__csr_io_decode_0_write_flush ; 
    wire core_id_illegal_insn =~ core_id_ctrl_legal |( core_id_ctrl_mul | core_id_ctrl_div )&~( core__csr_io_status_isa [12])| core_id_ctrl_amo &~( core__csr_io_status_isa [0])| core_id_ctrl_fp | core_id_ctrl_dp &~( core__csr_io_status_isa [3])| core__ibuf_io_inst_0_bits_rvc &~( core__csr_io_status_isa [2])| core_id_ctrl_rocc | core_id_csr_en &( core__csr_io_decode_0_read_illegal |~ core_id_csr_ren & core__csr_io_decode_0_write_illegal )|~ core__ibuf_io_inst_0_bits_rvc & core_id_system_insn & core__csr_io_decode_0_system_illegal ; 
    wire core_id_virtual_insn = core_id_ctrl_legal &( core_id_csr_en &~(~ core_id_csr_ren & core__csr_io_decode_0_write_illegal )& core__csr_io_decode_0_virtual_access_illegal |~ core__ibuf_io_inst_0_bits_rvc & core_id_system_insn & core__csr_io_decode_0_virtual_system_illegal ); 
    wire core_id_amo_aq = core__ibuf_io_inst_0_bits_inst_bits [26]; 
    wire core_id_amo_rl = core__ibuf_io_inst_0_bits_inst_bits [25]; 
    wire[3:0] core_id_fence_pred = core__ibuf_io_inst_0_bits_inst_bits [27:24]; 
    wire[3:0] core_id_fence_succ = core__ibuf_io_inst_0_bits_inst_bits [23:20]; 
    wire core_id_fence_next = core_id_ctrl_fence | core_id_ctrl_amo & core_id_amo_aq ; 
    wire core_id_mem_busy =~ core_io_dmem_ordered | core__io_dmem_req_valid_output ; 
    wire core_replay_wb_rocc = core_wb_reg_valid & core_wb_ctrl_rocc ; 
    wire core_id_do_fence = core_id_mem_busy &( core_id_ctrl_amo & core_id_amo_rl | core_id_ctrl_fence_i | core_id_reg_fence &( core_id_ctrl_mem | core_id_ctrl_rocc )); 
    wire core_id_xcpt = core__csr_io_interrupt | core__bpu_io_debug_if | core__bpu_io_xcpt_if | core__ibuf_io_inst_0_bits_xcpt0_pf_inst | core__ibuf_io_inst_0_bits_xcpt0_gf_inst | core__ibuf_io_inst_0_bits_xcpt0_ae_inst | core__ibuf_io_inst_0_bits_xcpt1_pf_inst | core__ibuf_io_inst_0_bits_xcpt1_gf_inst | core__ibuf_io_inst_0_bits_xcpt1_ae_inst | core_id_virtual_insn | core_id_illegal_insn ; 
    wire[31:0] core_id_cause = core__csr_io_interrupt  ?  core__csr_io_interrupt_cause :{27'h0, core__bpu_io_debug_if  ? 5'hE: core__bpu_io_xcpt_if  ? 5'h3: core__ibuf_io_inst_0_bits_xcpt0_pf_inst  ? 5'hC: core__ibuf_io_inst_0_bits_xcpt0_gf_inst  ? 5'h14: core__ibuf_io_inst_0_bits_xcpt0_ae_inst  ? 5'h1: core__ibuf_io_inst_0_bits_xcpt1_pf_inst  ? 5'hC: core__ibuf_io_inst_0_bits_xcpt1_gf_inst  ? 5'h14: core__ibuf_io_inst_0_bits_xcpt1_ae_inst  ? 5'h1: core_id_virtual_insn  ? 5'h16:5'h2}; 
    wire[4:0] core_ex_waddr = core_ex_reg_inst [11:7]; 
    wire[4:0] core_mem_waddr = core_mem_reg_inst [11:7]; 
    wire[4:0] core_wb_waddr = core_wb_reg_inst [11:7]; 
    wire[4:0] core_coreMonitorBundle_wrdst = core_wb_waddr ; 
    wire core__GEN_11 = core_ex_reg_valid & core_ex_ctrl_wxd ; 
    wire core__dcache_kill_mem_T = core_mem_reg_valid & core_mem_ctrl_wxd ; 
    wire core__GEN_12 = core__dcache_kill_mem_T &~ core_mem_ctrl_mem ; 
    wire core_id_bypass_src_0_0 =~(| core_id_raddr1 ); 
    wire core_id_bypass_src_0_1 = core__GEN_11 & core_ex_waddr == core_id_raddr1 ; 
    wire core__id_bypass_src_T_3 = core_mem_waddr == core_id_raddr1 ; 
    wire core_id_bypass_src_0_2 = core__GEN_12 & core__id_bypass_src_T_3 ; 
    wire core_id_bypass_src_0_3 = core__dcache_kill_mem_T & core__id_bypass_src_T_3 ; 
    wire core_id_bypass_src_1_0 =~(| core_id_raddr2 ); 
    wire core_id_bypass_src_1_1 = core__GEN_11 & core_ex_waddr == core_id_raddr2 ; 
    wire core__id_bypass_src_T_7 = core_mem_waddr == core_id_raddr2 ; 
    wire core_id_bypass_src_1_2 = core__GEN_12 & core__id_bypass_src_T_7 ; 
    wire core_id_bypass_src_1_3 = core__dcache_kill_mem_T & core__id_bypass_src_T_7 ; 
    reg core_ex_reg_rs_bypass_0 ; 
    reg core_ex_reg_rs_bypass_1 ; reg[1:0] core_ex_reg_rs_lsb_0 ; reg[1:0] core_ex_reg_rs_lsb_1 ; reg[29:0] core_ex_reg_rs_msb_0 ; reg[29:0] core_ex_reg_rs_msb_1 ; reg[31:0] core_casez_tmp ; 
  always @(*)
         begin 
             casez ( core_ex_reg_rs_lsb_0 )
              2 'b00: 
                  core_casez_tmp  =32'h0;
              2 'b01: 
                  core_casez_tmp  = core_mem_reg_wdata ;
              2 'b10: 
                  core_casez_tmp  = core_wb_reg_wdata ;
              default : 
                  core_casez_tmp  = core_dcache_bypass_data ;endcase
         end
    wire[31:0] core_ex_rs_0 = core_ex_reg_rs_bypass_0  ?  core_casez_tmp :{ core_ex_reg_rs_msb_0 , core_ex_reg_rs_lsb_0 }; reg[31:0] core_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( core_ex_reg_rs_lsb_1 )
              2 'b00: 
                  core_casez_tmp_0  =32'h0;
              2 'b01: 
                  core_casez_tmp_0  = core_mem_reg_wdata ;
              2 'b10: 
                  core_casez_tmp_0  = core_wb_reg_wdata ;
              default : 
                  core_casez_tmp_0  = core_dcache_bypass_data ;endcase
         end
    wire[31:0] core_ex_rs_1 = core_ex_reg_rs_bypass_1  ?  core_casez_tmp_0 :{ core_ex_reg_rs_msb_1 , core_ex_reg_rs_lsb_1 }; 
    wire core__ex_imm_b0_T_4 = core_ex_ctrl_sel_imm ==3'h5; 
    wire core_ex_imm_sign =~ core__ex_imm_b0_T_4 & core_ex_reg_inst [31]; 
    wire core_ex_imm_hi_hi_hi = core_ex_imm_sign ; 
    wire core__ex_imm_b4_1_T = core_ex_ctrl_sel_imm ==3'h2; 
    wire[10:0] core_ex_imm_b30_20 = core__ex_imm_b4_1_T  ?  core_ex_reg_inst [30:20]:{11{ core_ex_imm_sign }}; 
    wire[10:0] core_ex_imm_hi_hi_lo = core_ex_imm_b30_20 ; 
    wire[7:0] core_ex_imm_b19_12 = core_ex_ctrl_sel_imm !=3'h2& core_ex_ctrl_sel_imm !=3'h3 ? {8{ core_ex_imm_sign }}: core_ex_reg_inst [19:12]; 
    wire[7:0] core_ex_imm_hi_lo_hi = core_ex_imm_b19_12 ; 
    wire core__ex_imm_b4_1_T_2 = core_ex_ctrl_sel_imm ==3'h1; 
    wire core_ex_imm_b11 =~( core__ex_imm_b4_1_T | core__ex_imm_b0_T_4 )&( core_ex_ctrl_sel_imm ==3'h3 ?  core_ex_reg_inst [20]: core__ex_imm_b4_1_T_2  ?  core_ex_reg_inst [7]: core_ex_imm_sign ); 
    wire core_ex_imm_hi_lo_lo = core_ex_imm_b11 ; 
    wire[5:0] core_ex_imm_b10_5 = core__ex_imm_b4_1_T | core__ex_imm_b0_T_4  ? 6'h0: core_ex_reg_inst [30:25]; 
    wire core__ex_imm_b0_T = core_ex_ctrl_sel_imm ==3'h0; 
    wire[3:0] core_ex_imm_b4_1 = core__ex_imm_b4_1_T  ? 4'h0: core__ex_imm_b0_T | core__ex_imm_b4_1_T_2  ?  core_ex_reg_inst [11:8]: core__ex_imm_b0_T_4  ?  core_ex_reg_inst [19:16]: core_ex_reg_inst [24:21]; 
    wire core_ex_imm_b0 = core__ex_imm_b0_T  ?  core_ex_reg_inst [7]: core_ex_ctrl_sel_imm ==3'h4 ?  core_ex_reg_inst [20]: core__ex_imm_b0_T_4 & core_ex_reg_inst [15]; 
    wire[9:0] core_ex_imm_lo_hi ={ core_ex_imm_b10_5 , core_ex_imm_b4_1 }; 
    wire[10:0] core_ex_imm_lo ={ core_ex_imm_lo_hi , core_ex_imm_b0 }; 
    wire[8:0] core_ex_imm_hi_lo ={ core_ex_imm_hi_lo_hi , core_ex_imm_hi_lo_lo }; 
    wire[11:0] core_ex_imm_hi_hi ={ core_ex_imm_hi_hi_hi , core_ex_imm_hi_hi_lo }; 
    wire[20:0] core_ex_imm_hi ={ core_ex_imm_hi_hi , core_ex_imm_hi_lo }; 
    wire[31:0] core_ex_imm ={ core_ex_imm_hi , core_ex_imm_lo }; 
    wire[31:0] core_ex_op1 = core_ex_ctrl_sel_alu1 ==2'h2 ?  core_ex_reg_pc : core_ex_ctrl_sel_alu1 ==2'h1 ?  core_ex_rs_0 :32'h0; reg[31:0] core_casez_tmp_1 ; 
    wire[3:0] core__ex_op2_T_1 = core_ex_reg_rvc  ? 4'h2:4'h4; 
  always @(*)
         begin 
             casez ( core_ex_ctrl_sel_alu2 )
              2 'b00: 
                  core_casez_tmp_1  =32'h0;
              2 'b01: 
                  core_casez_tmp_1  ={{28{ core__ex_op2_T_1 [3]}}, core__ex_op2_T_1 };
              2 'b10: 
                  core_casez_tmp_1  = core_ex_rs_1 ;
              default : 
                  core_casez_tmp_1  = core_ex_imm ;endcase
         end
    wire[31:0] core_ex_op2 = core_casez_tmp_1 ; 
    wire core__div_io_req_valid_T = core_ex_reg_valid & core_ex_ctrl_div ; 
    wire[1:0] core_hi ={ core__ibuf_io_inst_0_bits_xcpt1_pf_inst , core__ibuf_io_inst_0_bits_xcpt1_gf_inst }; 
    wire[1:0] core_hi_1 ={ core__ibuf_io_inst_0_bits_xcpt0_pf_inst , core__ibuf_io_inst_0_bits_xcpt0_gf_inst }; 
    wire core_do_bypass = core_id_bypass_src_0_0 | core_id_bypass_src_0_1 | core_id_bypass_src_0_2 | core_id_bypass_src_0_3 ; 
    wire[1:0] core_bypass_src = core_id_bypass_src_0_0  ? 2'h0: core_id_bypass_src_0_1  ? 2'h1:{1'h1,~ core_id_bypass_src_0_2 }; 
    wire core_do_bypass_1 = core_id_bypass_src_1_0 | core_id_bypass_src_1_1 | core_id_bypass_src_1_2 | core_id_bypass_src_1_3 ; 
    wire[1:0] core_bypass_src_1 = core_id_bypass_src_1_0  ? 2'h0: core_id_bypass_src_1_1  ? 2'h1:{1'h1,~ core_id_bypass_src_1_2 }; 
    wire[31:0] core_inst = core__ibuf_io_inst_0_bits_rvc  ? {16'h0, core__ibuf_io_inst_0_bits_raw [15:0]}: core__ibuf_io_inst_0_bits_raw ; 
    wire core_ex_pc_valid = core_ex_reg_valid | core_ex_reg_replay | core_ex_reg_xcpt_interrupt ; 
    wire core_wb_dcache_miss = core_wb_ctrl_mem &~ core_io_dmem_resp_valid ; 
    wire core_replay_ex_structural = core_ex_ctrl_mem &~ core_io_dmem_req_ready | core_ex_ctrl_div &~ core__div_io_req_ready ; 
    wire core_replay_ex_load_use = core_wb_dcache_miss & core_ex_reg_load_use ; 
    wire core_replay_ex = core_ex_reg_replay | core_ex_reg_valid &( core_replay_ex_structural | core_replay_ex_load_use ); 
    wire core_ctrl_killx = core_take_pc_mem_wb | core_replay_ex |~ core_ex_reg_valid ; 
    wire core__mem_reg_store_T_3 = core_ex_ctrl_mem_cmd ==5'h7; 
    wire core_ex_slow_bypass = core__mem_reg_store_T_3 |~( core_ex_reg_mem_size [1]); 
    wire core_ex_xcpt = core_ex_reg_xcpt_interrupt | core_ex_reg_xcpt ; 
    wire core_mem_pc_valid = core_mem_reg_valid | core_mem_reg_replay | core_mem_reg_xcpt_interrupt ; 
    wire core__mem_cfi_taken_T = core_mem_ctrl_branch & core_mem_br_taken ; 
    wire core_mem_br_target_sign = core_mem_reg_inst [31]; 
    wire core_mem_br_target_sign_1 = core_mem_reg_inst [31]; 
    wire core_mem_br_target_hi_hi_hi = core_mem_br_target_sign ; 
    wire[10:0] core_mem_br_target_b30_20 ={11{ core_mem_br_target_sign }}; 
    wire[10:0] core_mem_br_target_hi_hi_lo = core_mem_br_target_b30_20 ; 
    wire[7:0] core_mem_br_target_b19_12_1 = core_mem_reg_inst [19:12]; 
    wire[7:0] core_mem_br_target_b19_12 ={8{ core_mem_br_target_sign }}; 
    wire[7:0] core_mem_br_target_hi_lo_hi = core_mem_br_target_b19_12 ; 
    wire core_mem_br_target_b11_1 = core_mem_reg_inst [20]; 
    wire core_mem_br_target_b11 = core_mem_reg_inst [7]; 
    wire core_mem_br_target_hi_lo_lo = core_mem_br_target_b11 ; 
    wire[5:0] core_mem_br_target_b10_5 = core_mem_reg_inst [30:25]; 
    wire[5:0] core_mem_br_target_b10_5_1 = core_mem_reg_inst [30:25]; 
    wire[3:0] core_mem_br_target_b4_1 = core_mem_reg_inst [11:8]; 
    wire[3:0] core_mem_br_target_b4_1_1 = core_mem_reg_inst [24:21]; 
    wire[9:0] core_mem_br_target_lo_hi ={ core_mem_br_target_b10_5 , core_mem_br_target_b4_1 }; 
    wire[10:0] core_mem_br_target_lo ={ core_mem_br_target_lo_hi ,1'h0}; 
    wire[8:0] core_mem_br_target_hi_lo ={ core_mem_br_target_hi_lo_hi , core_mem_br_target_hi_lo_lo }; 
    wire[11:0] core_mem_br_target_hi_hi ={ core_mem_br_target_hi_hi_hi , core_mem_br_target_hi_hi_lo }; 
    wire[20:0] core_mem_br_target_hi ={ core_mem_br_target_hi_hi , core_mem_br_target_hi_lo }; 
    wire core_mem_br_target_hi_hi_hi_1 = core_mem_br_target_sign_1 ; 
    wire[10:0] core_mem_br_target_b30_20_1 ={11{ core_mem_br_target_sign_1 }}; 
    wire[10:0] core_mem_br_target_hi_hi_lo_1 = core_mem_br_target_b30_20_1 ; 
    wire[7:0] core_mem_br_target_hi_lo_hi_1 = core_mem_br_target_b19_12_1 ; 
    wire core_mem_br_target_hi_lo_lo_1 = core_mem_br_target_b11_1 ; 
    wire[9:0] core_mem_br_target_lo_hi_1 ={ core_mem_br_target_b10_5_1 , core_mem_br_target_b4_1_1 }; 
    wire[10:0] core_mem_br_target_lo_1 ={ core_mem_br_target_lo_hi_1 ,1'h0}; 
    wire[8:0] core_mem_br_target_hi_lo_1 ={ core_mem_br_target_hi_lo_hi_1 , core_mem_br_target_hi_lo_lo_1 }; 
    wire[11:0] core_mem_br_target_hi_hi_1 ={ core_mem_br_target_hi_hi_hi_1 , core_mem_br_target_hi_hi_lo_1 }; 
    wire[20:0] core_mem_br_target_hi_1 ={ core_mem_br_target_hi_hi_1 , core_mem_br_target_hi_lo_1 }; 
    wire[3:0] core__mem_br_target_T_6 = core_mem_reg_rvc  ? 4'h2:4'h4; 
    wire[31:0] core_mem_br_target = core_mem_reg_pc +( core__mem_cfi_taken_T  ? { core_mem_br_target_hi , core_mem_br_target_lo }: core_mem_ctrl_jal  ? { core_mem_br_target_hi_1 , core_mem_br_target_lo_1 }:{{28{ core__mem_br_target_T_6 [3]}}, core__mem_br_target_T_6 }); 
    wire[31:0] core_mem_npc =( core_mem_ctrl_jalr  ?  core_mem_reg_wdata : core_mem_br_target )&32'hFFFFFFFE; 
    wire core_mem_wrong_npc = core_ex_pc_valid  ?  core_mem_npc != core_ex_reg_pc :~( core__ibuf_io_inst_0_valid | core_io_imem_resp_valid )| core_mem_npc != core__ibuf_io_pc ; 
    wire core_mem_npc_misaligned =~( core__csr_io_status_isa [2])& core_mem_npc [1]; 
    wire[31:0] core_mem_int_wdata =~ core_mem_reg_xcpt &( core_mem_ctrl_jalr ^ core_mem_npc_misaligned ) ?  core_mem_br_target : core_mem_reg_wdata ; 
    wire core_mem_cfi = core_mem_ctrl_branch | core_mem_ctrl_jalr | core_mem_ctrl_jal ; 
    wire core_mem_cfi_taken = core__mem_cfi_taken_T | core_mem_ctrl_jalr | core_mem_ctrl_jal ; 
    wire core_mem_direction_misprediction = core_mem_ctrl_branch & core_mem_br_taken ; 
  assign  core_take_pc_mem = core_mem_reg_valid &~ core_mem_reg_xcpt & core_mem_cfi_taken ; 
    wire[1:0] core_size = core_ex_ctrl_rocc  ? 2'h2: core_ex_reg_mem_size ; 
    wire[1:0] core_mem_reg_rs2_size = core_size ; 
    wire core_mem_breakpoint = core_mem_reg_load & core__bpu_io_xcpt_ld | core_mem_reg_store & core__bpu_io_xcpt_st ; 
    wire core_mem_debug_breakpoint = core_mem_reg_load & core__bpu_io_debug_ld | core_mem_reg_store & core__bpu_io_debug_st ; 
    wire core_mem_ldst_xcpt = core_mem_debug_breakpoint | core_mem_breakpoint ; 
    wire[3:0] core_mem_ldst_cause = core_mem_debug_breakpoint  ? 4'hE:4'h3; 
    wire core__GEN_13 = core_mem_reg_xcpt_interrupt | core_mem_reg_xcpt ; 
    wire core__GEN_14 = core_mem_reg_valid & core_mem_npc_misaligned ; 
    wire core_mem_xcpt = core__GEN_13 | core__GEN_14 | core_mem_reg_valid & core_mem_ldst_xcpt ; 
    wire[31:0] core_mem_cause = core__GEN_13  ?  core_mem_reg_cause :{28'h0, core__GEN_14  ? 4'h0: core_mem_ldst_cause }; 
    wire core_dcache_kill_mem = core__dcache_kill_mem_T & core_io_dmem_replay_next ; 
    wire core_replay_mem = core_dcache_kill_mem | core_mem_reg_replay ; 
    wire core_killm_common = core_dcache_kill_mem | core_take_pc_wb | core_mem_reg_xcpt |~ core_mem_reg_valid ; 
    reg core_div_io_kill_REG ; 
    wire core_ctrl_killm = core_killm_common | core_mem_xcpt ; 
    wire core__GEN_15 = core_wb_reg_valid & core_wb_ctrl_mem ; 
    wire core__GEN_16 = core__GEN_15 & core_io_dmem_s2_xcpt_pf_st ; 
    wire core__GEN_17 = core__GEN_15 & core_io_dmem_s2_xcpt_pf_ld ; 
    wire core__GEN_18 = core__GEN_15 & core_io_dmem_s2_xcpt_ae_st ; 
    wire core__GEN_19 = core__GEN_15 & core_io_dmem_s2_xcpt_ae_ld ; 
    wire core__GEN_20 = core__GEN_15 & core_io_dmem_s2_xcpt_ma_st ; 
    wire core_wb_xcpt = core_wb_reg_xcpt | core__GEN_16 | core__GEN_17 | core__GEN_18 | core__GEN_19 | core__GEN_20 | core__GEN_15 & core_io_dmem_s2_xcpt_ma_ld ; 
    wire[31:0] core_wb_cause = core_wb_reg_xcpt  ?  core_wb_reg_cause :{27'h0, core__GEN_16  ? 5'hF: core__GEN_17  ? 5'hD:{2'h0, core__GEN_18  ? 3'h7: core__GEN_19  ? 3'h5:{1'h1, core__GEN_20 ,1'h0}}}; 
    wire core_wb_pc_valid = core_wb_reg_valid | core_wb_reg_replay | core_wb_reg_xcpt ; 
    wire core_wb_wxd = core_wb_reg_valid & core_wb_ctrl_wxd ; 
    wire core_wb_set_sboard = core_wb_ctrl_div | core_wb_dcache_miss | core_wb_ctrl_rocc ; 
    wire core_replay_wb_common = core_io_dmem_s2_nack | core_wb_reg_replay ; 
    wire core_replay_wb = core_replay_wb_common | core_replay_wb_rocc ; 
  assign  core_take_pc_wb = core_replay_wb | core_wb_xcpt | core__csr_io_eret | core_wb_reg_flush_pipe ; 
    wire core_dmem_resp_fpu = core_io_dmem_resp_bits_tag [0]; 
    wire core_dmem_resp_xpu =~ core_dmem_resp_fpu ; 
    wire[4:0] core_dmem_resp_waddr = core_io_dmem_resp_bits_tag [5:1]; 
    wire core_dmem_resp_valid = core_io_dmem_resp_valid & core_io_dmem_resp_bits_has_data ; 
    wire core_dmem_resp_replay = core_dmem_resp_valid & core_io_dmem_resp_bits_replay ; 
    wire core__GEN_21 = core_dmem_resp_replay & core_dmem_resp_xpu ; 
  assign  core__GEN =~ core__GEN_21 &~ core_wb_wxd ; 
    wire[4:0] core_ll_waddr = core__GEN_21  ?  core_dmem_resp_waddr : core__div_io_resp_bits_tag ; 
    wire core_ll_wen = core__GEN_21 | core__GEN & core__div_io_resp_valid ; 
    wire core_wb_valid = core_wb_reg_valid &~ core_replay_wb &~ core_wb_xcpt ; 
    wire core_wb_wen = core_wb_valid & core_wb_ctrl_wxd ; 
    wire core_rf_wen = core_wb_wen | core_ll_wen ; 
    wire[4:0] core_rf_waddr = core_ll_wen  ?  core_ll_waddr : core_wb_waddr ; 
    wire[4:0] core_xrfWriteBundle_wrdst = core_rf_waddr ; 
    wire[31:0] core_ll_wdata ; 
    wire[31:0] core_rf_wdata = core_dmem_resp_valid & core_dmem_resp_xpu  ?  core_io_dmem_resp_bits_data : core_ll_wen  ?  core_ll_wdata :(| core_wb_ctrl_csr ) ?  core__csr_io_rw_rdata : core_wb_reg_wdata ; 
    wire[31:0] core_coreMonitorBundle_wrdata = core_rf_wdata ; 
    wire[31:0] core_xrfWriteBundle_wrdata = core_rf_wdata ; 
    wire[31:0] core_id_rs_0 = core_rf_wen &(| core_rf_waddr )& core_rf_waddr == core_id_raddr1  ?  core_rf_wdata : core__rf_ext_R1_data ; 
    wire[31:0] core_id_rs_1 = core_rf_wen &(| core_rf_waddr )& core_rf_waddr == core_id_raddr2  ?  core_rf_wdata : core__rf_ext_R0_data ; 
    wire core_tval_dmem_addr =~ core_wb_reg_xcpt ; 
    wire core__csr_io_htval_htval_valid_imem_T = core_wb_reg_cause ==32'h14; 
    wire core_tval_any_addr = core_tval_dmem_addr | core_wb_reg_cause ==32'h3| core_wb_reg_cause ==32'h1| core_wb_reg_cause ==32'hC| core__csr_io_htval_htval_valid_imem_T ; 
    wire core_tval_inst = core_wb_reg_cause ==32'h2; 
    wire core_tval_valid = core_wb_xcpt &( core_tval_any_addr | core_tval_inst ); 
    wire core_csr_io_htval_htval_valid_imem = core_wb_reg_xcpt & core__csr_io_htval_htval_valid_imem_T ; 
    wire[31:0] core_csr_io_htval_htval_imem = core_csr_io_htval_htval_valid_imem  ?  core_io_imem_gpa_bits :32'h0; 
    wire core__GEN_22 = core_id_ctrl_rxs1 &(| core_id_raddr1 ); 
    wire core__GEN_23 = core_id_ctrl_rxs2 &(| core_id_raddr2 ); 
    wire[4:0] core_id_waddr ; 
    wire core__GEN_24 = core_id_ctrl_wxd &(| core_id_waddr ); reg[31:0] core__r ; 
    wire[31:0] core_r ={ core__r [31:1],1'h0}; 
    wire[31:0] core__id_sboard_hazard_T = core_r >> core_id_raddr1 ; 
    wire[31:0] core__id_sboard_hazard_T_7 = core_r >> core_id_raddr2 ; 
    wire[31:0] core__id_sboard_hazard_T_14 = core_r >> core_id_waddr ; 
    wire core_id_sboard_hazard = core__GEN_22 & core__id_sboard_hazard_T [0]&~( core_ll_wen & core_ll_waddr == core_id_raddr1 )| core__GEN_23 & core__id_sboard_hazard_T_7 [0]&~( core_ll_wen & core_ll_waddr == core_id_raddr2 )| core__GEN_24 & core__id_sboard_hazard_T_14 [0]&~( core_ll_wen & core_ll_waddr == core_id_waddr ); 
    wire core_ex_cannot_bypass =(| core_ex_ctrl_csr )| core_ex_ctrl_jalr | core_ex_ctrl_mem | core_ex_ctrl_mul | core_ex_ctrl_div | core_ex_ctrl_fp | core_ex_ctrl_rocc ; 
    wire core_data_hazard_ex = core_ex_ctrl_wxd &( core__GEN_22 & core_id_raddr1 == core_ex_waddr | core__GEN_23 & core_id_raddr2 == core_ex_waddr | core__GEN_24 & core_id_waddr == core_ex_waddr ); 
    wire core_id_ex_hazard = core_ex_reg_valid & core_data_hazard_ex & core_ex_cannot_bypass ; 
    wire core_mem_cannot_bypass =(| core_mem_ctrl_csr )| core_mem_ctrl_mem & core_mem_mem_cmd_bh | core_mem_ctrl_mul | core_mem_ctrl_div | core_mem_ctrl_fp | core_mem_ctrl_rocc ; 
    wire core_data_hazard_mem = core_mem_ctrl_wxd &( core__GEN_22 & core_id_raddr1 == core_mem_waddr | core__GEN_23 & core_id_raddr2 == core_mem_waddr | core__GEN_24 & core_id_waddr == core_mem_waddr ); 
    wire core_id_mem_hazard = core_mem_reg_valid & core_data_hazard_mem & core_mem_cannot_bypass ; 
    wire core_id_load_use = core_mem_reg_valid & core_data_hazard_mem & core_mem_ctrl_mem ; 
    wire core_data_hazard_wb = core_wb_ctrl_wxd &( core__GEN_22 & core_id_raddr1 == core_wb_waddr | core__GEN_23 & core_id_raddr2 == core_wb_waddr | core__GEN_24 & core_id_waddr == core_wb_waddr ); 
    wire core_id_wb_hazard = core_wb_reg_valid & core_data_hazard_wb & core_wb_set_sboard ; 
    reg core_dcache_blocked_blocked ; 
    wire core_dcache_blocked = core_dcache_blocked_blocked &~ core_io_dmem_perf_grant ; 
    reg core_rocc_blocked ; 
    wire core_ctrl_stalld = core_id_ex_hazard | core_id_mem_hazard | core_id_wb_hazard | core_id_sboard_hazard | core__csr_io_singleStep &( core_ex_reg_valid | core_mem_reg_valid | core_wb_reg_valid )| core_id_ctrl_mem & core_dcache_blocked | core_id_ctrl_rocc & core_rocc_blocked | core_id_ctrl_div &(~( core__div_io_req_ready | core__div_io_resp_valid &~ core_wb_wxd )| core__div_io_req_valid_T )| core_id_do_fence | core__csr_io_csr_stall | core_id_reg_pause ; 
    wire core_ctrl_killd =~ core__ibuf_io_inst_0_valid | core__ibuf_io_inst_0_bits_replay | core_take_pc_mem_wb | core_ctrl_stalld | core__csr_io_interrupt ; 
    reg core_io_imem_progress_REG ; 
    wire core__io_imem_sfence_valid_output = core_wb_reg_valid & core_wb_reg_sfence ; 
  assign  core__io_dmem_req_valid_output = core_ex_reg_valid & core_ex_ctrl_mem ; 
    wire[5:0] core_ex_dcache_tag ={ core_ex_waddr , core_ex_ctrl_fp }; 
    wire core_unpause = core__csr_io_time [4:0]==5'h0| core__csr_io_inhibit_cycle | core_take_pc_mem_wb ; 
    reg core_icache_blocked_REG ; 
    wire core_icache_blocked =~( core_io_imem_resp_valid | core_icache_blocked_REG ); 
    wire[31:0] core__GEN_25 ={31'h0, core_io_hartid }; 
    wire[31:0] core_coreMonitorBundle_hartid ; 
  assign  core_coreMonitorBundle_hartid = core__GEN_25 ; 
    wire[31:0] core_xrfWriteBundle_hartid ; 
  assign  core_xrfWriteBundle_hartid = core__GEN_25 ; 
    wire core_coreMonitorBundle_valid = core__csr_io_trace_0_valid &~ core__csr_io_trace_0_exception ; 
    wire core_coreMonitorBundle_wrenx = core_wb_wen &~ core_wb_set_sboard ; 
    wire[4:0] core_coreMonitorBundle_rd0src = core_wb_reg_inst [19:15]; reg[31:0] core_coreMonitorBundle_rd0val_REG ; reg[31:0] core_coreMonitorBundle_rd0val_REG_1 ; 
    wire[31:0] core_coreMonitorBundle_rd0val = core_coreMonitorBundle_rd0val_REG_1 ; 
    wire[4:0] core_coreMonitorBundle_rd1src = core_wb_reg_inst [24:20]; reg[31:0] core_coreMonitorBundle_rd1val_REG ; reg[31:0] core_coreMonitorBundle_rd1val_REG_1 ; 
    wire[31:0] core_coreMonitorBundle_timer ; 
    wire[31:0] core_coreMonitorBundle_pc ; 
    wire[31:0] core_coreMonitorBundle_rd1val = core_coreMonitorBundle_rd1val_REG_1 ; 
    wire[31:0] core_coreMonitorBundle_inst ; 
    wire core__GEN_26 = core_wb_ctrl_rxs1 | core_wb_ctrl_rfs1 ; 
    wire core__GEN_27 = core_wb_ctrl_rxs2 | core_wb_ctrl_rfs2 ; 
  always @( posedge  core_clock )
         begin 
             if (~ core_reset &~(~ core_csr_io_htval_htval_valid_imem | core_io_imem_gpa_valid ))
                 begin 
                     if (1)$error("Assertion failed\n    at RocketCore.scala:718 assert(!htval_valid_imem || io.imem.gpa.valid)\n");
                     if (1)$fatal;
                 end 
             if ((1)& core__csr_io_trace_0_valid &~ core_reset )$fwrite(32'h80000002,"C%d: %d [%d] pc=[%x] W[r%d=%x][%d] R[r%d=%x] R[r%d=%x] inst=[%x] DASM(%x)\n", core_io_hartid , core_coreMonitorBundle_timer , core_coreMonitorBundle_valid , core_coreMonitorBundle_pc , core_wb_ctrl_wxd | core_wb_ctrl_wfd  ?  core_coreMonitorBundle_wrdst :5'h0, core_coreMonitorBundle_wrenx  ?  core_coreMonitorBundle_wrdata :32'h0, core_coreMonitorBundle_wrenx , core__GEN_26  ?  core_coreMonitorBundle_rd0src :5'h0, core__GEN_26  ?  core_coreMonitorBundle_rd0val :32'h0, core__GEN_27  ?  core_coreMonitorBundle_rd1src :5'h0, core__GEN_27  ?  core_coreMonitorBundle_rd1val :32'h0, core_coreMonitorBundle_inst , core_coreMonitorBundle_inst );
         end
    wire core_xrfWriteBundle_wrenx = core_rf_wen &~( core__csr_io_trace_0_valid & core_wb_wen & core_wb_waddr == core_rf_waddr ); 
    wire[2:0] core__GEN_28 ={ core_hi , core__ibuf_io_inst_0_bits_xcpt1_ae_inst }; 
    wire core__GEN_29 = core__bpu_io_xcpt_if |(|{ core_hi_1 , core__ibuf_io_inst_0_bits_xcpt0_ae_inst }); 
    wire core__GEN_30 = core_id_ctrl_mem_cmd ==5'h14; 
    wire core__GEN_31 = core_id_ctrl_rxs1 &~ core_do_bypass ; 
    wire core__GEN_32 = core_id_illegal_insn | core_id_virtual_insn ; 
    wire core__mem_reg_store_T_5 = core_ex_ctrl_mem_cmd ==5'h4; 
    wire core__mem_reg_store_T_6 = core_ex_ctrl_mem_cmd ==5'h9; 
    wire core__mem_reg_store_T_7 = core_ex_ctrl_mem_cmd ==5'hA; 
    wire core__mem_reg_store_T_8 = core_ex_ctrl_mem_cmd ==5'hB; 
    wire core__mem_reg_store_T_12 = core_ex_ctrl_mem_cmd ==5'h8; 
    wire core__mem_reg_store_T_13 = core_ex_ctrl_mem_cmd ==5'hC; 
    wire core__mem_reg_store_T_14 = core_ex_ctrl_mem_cmd ==5'hD; 
    wire core__mem_reg_store_T_15 = core_ex_ctrl_mem_cmd ==5'hE; 
    wire core__mem_reg_store_T_16 = core_ex_ctrl_mem_cmd ==5'hF; 
    wire[31:0] core__GEN_33 = core_r &~( core_ll_wen  ? 32'h1<< core_ll_waddr :32'h0); 
    wire core__GEN_34 = core_wb_set_sboard & core_wb_wen ; 
    wire core__GEN_35 = core_id_ctrl_rxs2 &~ core_do_bypass_1 ; 
    wire core__GEN_36 = core_mem_reg_valid & core_mem_reg_flush_pipe ; 
    wire core__GEN_37 = core__GEN_36 |~ core_ex_pc_valid ; 
    wire core__GEN_38 = core_ex_ctrl_jalr & core__csr_io_status_debug ; 
  always @( posedge  core_clock )
         begin  
             core_id_reg_pause  <=~ core_unpause &(~ core_ctrl_killd & core_id_ctrl_fence & core_id_fence_succ ==4'h0| core_id_reg_pause ); 
             core_imem_might_request_reg  <= core_ex_pc_valid | core_mem_pc_valid | core__csr_io_customCSRs_0_value [1];
             if ( core_ctrl_killd )
                 begin 
                 end 
              else 
                 begin  
                     core_ex_ctrl_legal  <= core_id_ctrl_legal ; 
                     core_ex_ctrl_fp  <= core_id_ctrl_fp ; 
                     core_ex_ctrl_rocc  <= core_id_ctrl_rocc ; 
                     core_ex_ctrl_branch  <= core_id_ctrl_branch ; 
                     core_ex_ctrl_jal  <= core_id_ctrl_jal ; 
                     core_ex_ctrl_jalr  <= core_id_ctrl_jalr ; 
                     core_ex_ctrl_rxs2  <= core_id_ctrl_rxs2 ; 
                     core_ex_ctrl_rxs1  <= core_id_ctrl_rxs1 ; 
                     core_ex_ctrl_sel_alu2  <= core_id_xcpt  ? ( core__GEN_29  ? 2'h0:{1'h0,| core__GEN_28 }): core_id_ctrl_sel_alu2 ; 
                     core_ex_ctrl_sel_alu1  <= core_id_xcpt  ? ( core__GEN_29 |(| core__GEN_28 ) ? 2'h2:2'h1): core_id_ctrl_sel_alu1 ; 
                     core_ex_ctrl_sel_imm  <= core_id_ctrl_sel_imm ; 
                     core_ex_ctrl_alu_dw  <= core_id_xcpt | core_id_ctrl_alu_dw ; 
                     core_ex_ctrl_alu_fn  <= core_id_xcpt  ? 4'h0: core_id_ctrl_alu_fn ; 
                     core_ex_ctrl_mem  <= core_id_ctrl_mem ; 
                     core_ex_ctrl_mem_cmd  <= core__GEN_30 & core__csr_io_status_v  ? 5'h15: core_id_ctrl_mem_cmd ; 
                     core_ex_ctrl_rfs1  <= core_id_ctrl_rfs1 ; 
                     core_ex_ctrl_rfs2  <= core_id_ctrl_rfs2 ; 
                     core_ex_ctrl_rfs3  <= core_id_ctrl_rfs3 ; 
                     core_ex_ctrl_wfd  <= core_id_ctrl_wfd ; 
                     core_ex_ctrl_mul  <= core_id_ctrl_mul ; 
                     core_ex_ctrl_div  <= core_id_ctrl_div ; 
                     core_ex_ctrl_wxd  <= core_id_ctrl_wxd ; 
                     core_ex_ctrl_csr  <= core_id_csr ; 
                     core_ex_ctrl_fence_i  <= core_id_ctrl_fence_i ; 
                     core_ex_ctrl_fence  <= core_id_ctrl_fence ; 
                     core_ex_ctrl_amo  <= core_id_ctrl_amo ; 
                     core_ex_ctrl_dp  <= core_id_ctrl_dp ; 
                     core_ex_reg_rvc  <= core_id_xcpt &(| core__GEN_28 )| core__ibuf_io_inst_0_bits_rvc ; 
                     core_ex_reg_flush_pipe  <= core_id_ctrl_fence_i | core_id_csr_flush ; 
                     core_ex_reg_load_use  <= core_id_load_use ; 
                     core_ex_reg_mem_size  <= core__GEN_30 | core_id_ctrl_mem_cmd ==5'h15| core_id_ctrl_mem_cmd ==5'h16| core_id_ctrl_mem_cmd ==5'h5 ? {| core_id_raddr2 ,| core_id_raddr1 }: core__ibuf_io_inst_0_bits_inst_bits [13:12]; 
                     core_ex_reg_rs_bypass_0  <=~ core__GEN_32 & core_do_bypass ; 
                     core_ex_reg_rs_bypass_1  <= core_do_bypass_1 ; 
                     core_ex_reg_rs_lsb_0  <= core__GEN_32  ?  core_inst [1:0]: core__GEN_31  ?  core_id_rs_0 [1:0]: core_bypass_src ; 
                     core_ex_reg_rs_lsb_1  <= core__GEN_35  ?  core_id_rs_1 [1:0]: core_bypass_src_1 ;
                     if ( core__GEN_32 ) 
                         core_ex_reg_rs_msb_0  <= core_inst [31:2];
                      else 
                         if ( core__GEN_31 ) 
                             core_ex_reg_rs_msb_0  <= core_id_rs_0 [31:2];
                 end 
             if ( core__GEN_37 )
                 begin 
                 end 
              else 
                 begin  
                     core_mem_ctrl_legal  <= core_ex_ctrl_legal ; 
                     core_mem_ctrl_fp  <= core_ex_ctrl_fp ; 
                     core_mem_ctrl_rocc  <= core_ex_ctrl_rocc ; 
                     core_mem_ctrl_branch  <= core_ex_ctrl_branch ; 
                     core_mem_ctrl_jal  <= core_ex_ctrl_jal ; 
                     core_mem_ctrl_jalr  <= core_ex_ctrl_jalr ; 
                     core_mem_ctrl_rxs2  <= core_ex_ctrl_rxs2 ; 
                     core_mem_ctrl_rxs1  <= core_ex_ctrl_rxs1 ; 
                     core_mem_ctrl_sel_alu2  <= core_ex_ctrl_sel_alu2 ; 
                     core_mem_ctrl_sel_alu1  <= core_ex_ctrl_sel_alu1 ; 
                     core_mem_ctrl_sel_imm  <= core_ex_ctrl_sel_imm ; 
                     core_mem_ctrl_alu_dw  <= core_ex_ctrl_alu_dw ; 
                     core_mem_ctrl_alu_fn  <= core_ex_ctrl_alu_fn ; 
                     core_mem_ctrl_mem  <= core_ex_ctrl_mem ; 
                     core_mem_ctrl_mem_cmd  <= core_ex_ctrl_mem_cmd ; 
                     core_mem_ctrl_rfs1  <= core_ex_ctrl_rfs1 ; 
                     core_mem_ctrl_rfs2  <= core_ex_ctrl_rfs2 ; 
                     core_mem_ctrl_rfs3  <= core_ex_ctrl_rfs3 ; 
                     core_mem_ctrl_wfd  <= core_ex_ctrl_wfd ; 
                     core_mem_ctrl_mul  <= core_ex_ctrl_mul ; 
                     core_mem_ctrl_div  <= core_ex_ctrl_div ; 
                     core_mem_ctrl_wxd  <= core_ex_ctrl_wxd ; 
                     core_mem_ctrl_csr  <= core_ex_ctrl_csr ; 
                     core_mem_ctrl_fence_i  <= core__GEN_38 | core_ex_ctrl_fence_i ; 
                     core_mem_ctrl_fence  <= core_ex_ctrl_fence ; 
                     core_mem_ctrl_amo  <= core_ex_ctrl_amo ; 
                     core_mem_ctrl_dp  <= core_ex_ctrl_dp ;
                 end 
             if ( core_mem_pc_valid )
                 begin  
                     core_wb_ctrl_legal  <= core_mem_ctrl_legal ; 
                     core_wb_ctrl_fp  <= core_mem_ctrl_fp ; 
                     core_wb_ctrl_rocc  <= core_mem_ctrl_rocc ; 
                     core_wb_ctrl_branch  <= core_mem_ctrl_branch ; 
                     core_wb_ctrl_jal  <= core_mem_ctrl_jal ; 
                     core_wb_ctrl_jalr  <= core_mem_ctrl_jalr ; 
                     core_wb_ctrl_rxs2  <= core_mem_ctrl_rxs2 ; 
                     core_wb_ctrl_rxs1  <= core_mem_ctrl_rxs1 ; 
                     core_wb_ctrl_sel_alu2  <= core_mem_ctrl_sel_alu2 ; 
                     core_wb_ctrl_sel_alu1  <= core_mem_ctrl_sel_alu1 ; 
                     core_wb_ctrl_sel_imm  <= core_mem_ctrl_sel_imm ; 
                     core_wb_ctrl_alu_dw  <= core_mem_ctrl_alu_dw ; 
                     core_wb_ctrl_alu_fn  <= core_mem_ctrl_alu_fn ; 
                     core_wb_ctrl_mem  <= core_mem_ctrl_mem ; 
                     core_wb_ctrl_mem_cmd  <= core_mem_ctrl_mem_cmd ; 
                     core_wb_ctrl_rfs1  <= core_mem_ctrl_rfs1 ; 
                     core_wb_ctrl_rfs2  <= core_mem_ctrl_rfs2 ; 
                     core_wb_ctrl_rfs3  <= core_mem_ctrl_rfs3 ; 
                     core_wb_ctrl_wfd  <= core_mem_ctrl_wfd ; 
                     core_wb_ctrl_mul  <= core_mem_ctrl_mul ; 
                     core_wb_ctrl_div  <= core_mem_ctrl_div ; 
                     core_wb_ctrl_wxd  <= core_mem_ctrl_wxd ; 
                     core_wb_ctrl_csr  <= core_mem_ctrl_csr ; 
                     core_wb_ctrl_fence_i  <= core_mem_ctrl_fence_i ; 
                     core_wb_ctrl_fence  <= core_mem_ctrl_fence ; 
                     core_wb_ctrl_amo  <= core_mem_ctrl_amo ; 
                     core_wb_ctrl_dp  <= core_mem_ctrl_dp ; 
                     core_wb_reg_cause  <= core_mem_cause ; 
                     core_wb_reg_pc  <= core_mem_reg_pc ; 
                     core_wb_reg_mem_size  <= core_mem_reg_mem_size ; 
                     core_wb_reg_hls_or_dv  <= core_mem_reg_hls_or_dv ; 
                     core_wb_reg_hfence_v  <= core_mem_ctrl_mem_cmd ==5'h15; 
                     core_wb_reg_hfence_g  <= core_mem_ctrl_mem_cmd ==5'h16; 
                     core_wb_reg_inst  <= core_mem_reg_inst ; 
                     core_wb_reg_raw_inst  <= core_mem_reg_raw_inst ; 
                     core_wb_reg_wdata  <=~ core_mem_reg_xcpt & core_mem_ctrl_fp & core_mem_ctrl_wxd  ? 32'h0: core_mem_int_wdata ; 
                     core_wb_reg_wphit_0  <= core_mem_reg_wphit_0 | core__bpu_io_bpwatch_0_rvalid_0 & core_mem_reg_load | core__bpu_io_bpwatch_0_wvalid_0 & core_mem_reg_store ;
                 end  
             core_ex_reg_xcpt_interrupt  <=~ core_take_pc_mem_wb & core__ibuf_io_inst_0_valid & core__csr_io_interrupt ; 
             core_ex_reg_valid  <=~ core_ctrl_killd ;
             if (~ core_ctrl_killd | core__csr_io_interrupt | core__ibuf_io_inst_0_bits_replay )
                 begin  
                     core_ex_reg_btb_resp_cfiType  <= core__ibuf_io_btb_resp_cfiType ; 
                     core_ex_reg_btb_resp_taken  <= core__ibuf_io_btb_resp_taken ; 
                     core_ex_reg_btb_resp_mask  <= core__ibuf_io_btb_resp_mask ; 
                     core_ex_reg_btb_resp_bridx  <= core__ibuf_io_btb_resp_bridx ; 
                     core_ex_reg_btb_resp_target  <= core__ibuf_io_btb_resp_target ; 
                     core_ex_reg_btb_resp_entry  <= core__ibuf_io_btb_resp_entry ; 
                     core_ex_reg_btb_resp_bht_history  <= core__ibuf_io_btb_resp_bht_history ; 
                     core_ex_reg_btb_resp_bht_value  <= core__ibuf_io_btb_resp_bht_value ; 
                     core_ex_reg_cause  <= core_id_cause ; 
                     core_ex_reg_pc  <= core__ibuf_io_pc ; 
                     core_ex_reg_inst  <= core__ibuf_io_inst_0_bits_inst_bits ; 
                     core_ex_reg_raw_inst  <= core__ibuf_io_inst_0_bits_raw ; 
                     core_ex_reg_wphit_0  <= core__bpu_io_bpwatch_0_ivalid_0 ;
                 end  
             core_ex_reg_xcpt  <=~ core_ctrl_killd & core_id_xcpt ; 
             core_ex_reg_replay  <=~ core_take_pc_mem_wb & core__ibuf_io_inst_0_valid & core__ibuf_io_inst_0_bits_replay ; 
             core_mem_reg_xcpt_interrupt  <=~ core_take_pc_mem_wb & core_ex_reg_xcpt_interrupt ; 
             core_mem_reg_valid  <=~ core_ctrl_killx ;
             if ( core__GEN_37 )
                 begin 
                 end 
              else 
                 begin  
                     core_mem_reg_rvc  <= core_ex_reg_rvc ; 
                     core_mem_reg_btb_resp_cfiType  <= core_ex_reg_btb_resp_cfiType ; 
                     core_mem_reg_btb_resp_taken  <= core_ex_reg_btb_resp_taken ; 
                     core_mem_reg_btb_resp_mask  <= core_ex_reg_btb_resp_mask ; 
                     core_mem_reg_btb_resp_bridx  <= core_ex_reg_btb_resp_bridx ; 
                     core_mem_reg_btb_resp_target  <= core_ex_reg_btb_resp_target ; 
                     core_mem_reg_btb_resp_entry  <= core_ex_reg_btb_resp_entry ; 
                     core_mem_reg_btb_resp_bht_history  <= core_ex_reg_btb_resp_bht_history ; 
                     core_mem_reg_btb_resp_bht_value  <= core_ex_reg_btb_resp_bht_value ;
                 end  
             core_mem_reg_xcpt  <=~ core_ctrl_killx & core_ex_xcpt ; 
             core_mem_reg_replay  <=~ core_take_pc_mem_wb & core_replay_ex ;
             if ( core__GEN_37 )
                 begin 
                 end 
              else 
                 begin  
                     core_mem_reg_flush_pipe  <= core__GEN_38 | core_ex_reg_flush_pipe ; 
                     core_mem_reg_cause  <= core_ex_reg_cause ; 
                     core_mem_reg_slow_bypass  <= core_ex_slow_bypass ; 
                     core_mem_reg_load  <= core_ex_ctrl_mem &( core_ex_ctrl_mem_cmd ==5'h0| core_ex_ctrl_mem_cmd ==5'h10| core_ex_ctrl_mem_cmd ==5'h6| core__mem_reg_store_T_3 | core__mem_reg_store_T_5 | core__mem_reg_store_T_6 | core__mem_reg_store_T_7 | core__mem_reg_store_T_8 | core__mem_reg_store_T_12 | core__mem_reg_store_T_13 | core__mem_reg_store_T_14 | core__mem_reg_store_T_15 | core__mem_reg_store_T_16 ); 
                     core_mem_reg_store  <= core_ex_ctrl_mem &( core_ex_ctrl_mem_cmd ==5'h1| core_ex_ctrl_mem_cmd ==5'h11| core__mem_reg_store_T_3 | core__mem_reg_store_T_5 | core__mem_reg_store_T_6 | core__mem_reg_store_T_7 | core__mem_reg_store_T_8 | core__mem_reg_store_T_12 | core__mem_reg_store_T_13 | core__mem_reg_store_T_14 | core__mem_reg_store_T_15 | core__mem_reg_store_T_16 ); 
                     core_mem_reg_pc  <= core_ex_reg_pc ; 
                     core_mem_reg_inst  <= core_ex_reg_inst ; 
                     core_mem_reg_mem_size  <= core_ex_reg_mem_size ; 
                     core_mem_reg_hls_or_dv  <= core__csr_io_status_dv ; 
                     core_mem_reg_raw_inst  <= core_ex_reg_raw_inst ; 
                     core_mem_reg_wdata  <= core__alu_io_out ;
                 end 
             if ( core__GEN_36 |~( core_ex_pc_valid & core_ex_ctrl_rxs2 &( core_ex_ctrl_mem | core_ex_ctrl_rocc )))
                 begin 
                 end 
              else  
                 core_mem_reg_rs2  <= core_mem_reg_rs2_size ==2'h0 ? {2{{2{ core_ex_rs_1 [7:0]}}}}: core_mem_reg_rs2_size ==2'h1 ? {2{ core_ex_rs_1 [15:0]}}: core_ex_rs_1 ;
             if ( core__GEN_37 )
                 begin 
                 end 
              else 
                 begin  
                     core_mem_br_taken  <= core__alu_io_cmp_out ; 
                     core_mem_reg_wphit_0  <= core_ex_reg_wphit_0 ;
                 end  
             core_wb_reg_valid  <=~ core_ctrl_killm ; 
             core_wb_reg_xcpt  <= core_mem_xcpt &~ core_take_pc_wb ; 
             core_wb_reg_replay  <= core_replay_mem &~ core_take_pc_wb ; 
             core_wb_reg_flush_pipe  <=~ core_ctrl_killm & core_mem_reg_flush_pipe ; 
             core_wb_reg_sfence  <=~ core_mem_pc_valid & core_wb_reg_sfence ;
             if ( core_mem_pc_valid & core_mem_ctrl_rocc ) 
                 core_wb_reg_rs2  <= core_mem_reg_rs2 ;
             if (~ core_ctrl_killd & core__GEN_35 ) 
                 core_ex_reg_rs_msb_1  <= core_id_rs_1 [31:2]; 
             core_div_io_kill_REG  <= core__div_io_req_ready & core__div_io_req_valid_T ; 
             core_dcache_blocked_blocked  <=~ core_io_dmem_req_ready &~ core_io_dmem_perf_grant &( core_dcache_blocked_blocked | core__io_dmem_req_valid_output | core_io_dmem_s2_nack ); 
             core_rocc_blocked  <=~ core_wb_xcpt &( core_replay_wb_rocc &~ core_replay_wb_common | core_rocc_blocked ); 
             core_io_imem_progress_REG  <= core_wb_reg_valid &~ core_replay_wb_common ; 
             core_icache_blocked_REG  <= core_io_imem_resp_valid ; 
             core_coreMonitorBundle_rd0val_REG  <= core_ex_rs_0 ; 
             core_coreMonitorBundle_rd0val_REG_1  <= core_coreMonitorBundle_rd0val_REG ; 
             core_coreMonitorBundle_rd1val_REG  <= core_ex_rs_1 ; 
             core_coreMonitorBundle_rd1val_REG_1  <= core_coreMonitorBundle_rd1val_REG ;
             if ( core_reset )
                 begin  
                     core_id_reg_fence  <=1'h0; 
                     core__r  <=32'h0;
                 end 
              else 
                 begin  
                     core_id_reg_fence  <=~ core_ctrl_killd & core_id_fence_next | core_id_mem_busy & core_id_reg_fence ;
                     if ( core_ll_wen | core__GEN_34 ) 
                         core__r  <= core__GEN_33 |( core__GEN_34  ? 32'h1<< core_wb_waddr :32'h0);
                      else 
                         if ( core_ll_wen ) 
                             core__r  <= core__GEN_33 ;
                 end 
         end
    wire core_ibuf_clock;
    wire core_ibuf_reset;
    wire core_ibuf_io_imem_ready;
    wire core_ibuf_io_imem_valid;
    wire[1:0] core_ibuf_io_imem_bits_btb_cfiType;
    wire core_ibuf_io_imem_bits_btb_taken;
    wire[1:0] core_ibuf_io_imem_bits_btb_mask;
    wire core_ibuf_io_imem_bits_btb_bridx;
    wire[31:0] core_ibuf_io_imem_bits_btb_target;
    wire core_ibuf_io_imem_bits_btb_entry;
    wire[7:0] core_ibuf_io_imem_bits_btb_bht_history;
    wire core_ibuf_io_imem_bits_btb_bht_value;
    wire[31:0] core_ibuf_io_imem_bits_pc;
    wire[31:0] core_ibuf_io_imem_bits_data;
    wire[1:0] core_ibuf_io_imem_bits_mask;
    wire core_ibuf_io_imem_bits_xcpt_pf_inst;
    wire core_ibuf_io_imem_bits_xcpt_gf_inst;
    wire core_ibuf_io_imem_bits_xcpt_ae_inst;
    wire core_ibuf_io_imem_bits_replay;
    wire core_ibuf_io_kill;
    wire[31:0] core_ibuf_io_pc;
    wire[1:0] core_ibuf_io_btb_resp_cfiType;
    wire core_ibuf_io_btb_resp_taken;
    wire[1:0] core_ibuf_io_btb_resp_mask;
    wire core_ibuf_io_btb_resp_bridx;
    wire[31:0] core_ibuf_io_btb_resp_target;
    wire core_ibuf_io_btb_resp_entry;
    wire[7:0] core_ibuf_io_btb_resp_bht_history;
    wire core_ibuf_io_btb_resp_bht_value;
    wire core_ibuf_io_inst_0_ready;
    wire core_ibuf_io_inst_0_valid;
    wire core_ibuf_io_inst_0_bits_xcpt0_pf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt0_gf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt0_ae_inst;
    wire core_ibuf_io_inst_0_bits_xcpt1_pf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt1_gf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt1_ae_inst;
    wire core_ibuf_io_inst_0_bits_replay;
    wire core_ibuf_io_inst_0_bits_rvc;
    wire[31:0] core_ibuf_io_inst_0_bits_inst_bits;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rd;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rs1;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rs2;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rs3;
    wire[31:0] core_ibuf_io_inst_0_bits_raw;

    wire core_ibuf__exp_io_rvc ; 
    reg core_ibuf_nBufValid ; reg[1:0] core_ibuf_buf_btb_cfiType ; 
    reg core_ibuf_buf_btb_taken ; reg[1:0] core_ibuf_buf_btb_mask ; 
    reg core_ibuf_buf_btb_bridx ; reg[31:0] core_ibuf_buf_btb_target ; 
    reg core_ibuf_buf_btb_entry ; reg[7:0] core_ibuf_buf_btb_bht_history ; 
    reg core_ibuf_buf_btb_bht_value ; reg[31:0] core_ibuf_buf_pc ; reg[31:0] core_ibuf_buf_data ; reg[1:0] core_ibuf_buf_mask ; 
    reg core_ibuf_buf_xcpt_pf_inst ; 
    reg core_ibuf_buf_xcpt_gf_inst ; 
    reg core_ibuf_buf_xcpt_ae_inst ; 
    reg core_ibuf_buf_replay ; reg[1:0] core_ibuf_ibufBTBResp_cfiType ; 
    reg core_ibuf_ibufBTBResp_taken ; reg[1:0] core_ibuf_ibufBTBResp_mask ; 
    reg core_ibuf_ibufBTBResp_bridx ; reg[31:0] core_ibuf_ibufBTBResp_target ; 
    reg core_ibuf_ibufBTBResp_entry ; reg[7:0] core_ibuf_ibufBTBResp_bht_history ; 
    reg core_ibuf_ibufBTBResp_bht_value ; 
    wire core_ibuf_pcWordBits = core_ibuf_io_imem_bits_pc [1]; 
    wire[1:0] core_ibuf__GEN ={1'h0, core_ibuf_pcWordBits }; 
    wire[1:0] core_ibuf_nIC =( core_ibuf_io_imem_bits_btb_taken  ? {1'h0, core_ibuf_io_imem_bits_btb_bridx }+2'h1:2'h2)- core_ibuf__GEN ; 
    wire[1:0] core_ibuf__GEN_0 ={1'h0, core_ibuf_nBufValid }; 
    wire[1:0] core_ibuf_nReady ; 
    wire[1:0] core_ibuf_nICReady = core_ibuf_nReady - core_ibuf__GEN_0 ; 
    wire[1:0] core_ibuf_nValid =( core_ibuf_io_imem_valid  ?  core_ibuf_nIC :2'h0)+ core_ibuf__GEN_0 ; 
    wire core_ibuf__nBufValid_T = core_ibuf_nReady >= core_ibuf__GEN_0 ; 
    wire[1:0] core_ibuf__nBufValid_T_6 = core_ibuf_nIC - core_ibuf_nICReady ; 
    wire[1:0] core_ibuf_shamt = core_ibuf__GEN + core_ibuf_nICReady ; 
    wire[63:0] core_ibuf_buf_data_data ={{2{ core_ibuf_io_imem_bits_data [31:16]}}, core_ibuf_io_imem_bits_data }; 
    wire[1:0] core_ibuf_icShiftAmt = core_ibuf__GEN_0 -2'h2- core_ibuf__GEN ; 
    wire[127:0] core_ibuf_icData_data ={{2{{2{ core_ibuf_io_imem_bits_data [31:16]}}}}, core_ibuf_io_imem_bits_data ,{2{ core_ibuf_io_imem_bits_data [15:0]}}}; 
    wire[190:0] core_ibuf__icData_T_4 ={63'h0, core_ibuf_icData_data }<<{185'h0, core_ibuf_icShiftAmt ,4'h0}; 
    wire[31:0] core_ibuf_icData = core_ibuf__icData_T_4 [95:64]; 
    wire[62:0] core_ibuf__icMask_T_2 =63'hFFFFFFFF<<{58'h0, core_ibuf_nBufValid ,4'h0}; 
    wire[31:0] core_ibuf_icMask = core_ibuf__icMask_T_2 [31:0]; 
    wire[31:0] core_ibuf_inst = core_ibuf_icData & core_ibuf_icMask | core_ibuf_buf_data &~ core_ibuf_icMask ; 
    wire[3:0] core_ibuf__valid_T =4'h1<< core_ibuf_nValid ; 
    wire[1:0] core_ibuf_valid = core_ibuf__valid_T [1:0]-2'h1; 
    wire[1:0] core_ibuf_bufMask =(2'h1<< core_ibuf__GEN_0 )-2'h1; 
    wire core_ibuf_xcpt_0_pf_inst = core_ibuf_bufMask [0] ?  core_ibuf_buf_xcpt_pf_inst : core_ibuf_io_imem_bits_xcpt_pf_inst ; 
    wire core_ibuf_xcpt_0_gf_inst = core_ibuf_bufMask [0] ?  core_ibuf_buf_xcpt_gf_inst : core_ibuf_io_imem_bits_xcpt_gf_inst ; 
    wire core_ibuf_xcpt_0_ae_inst = core_ibuf_bufMask [0] ?  core_ibuf_buf_xcpt_ae_inst : core_ibuf_io_imem_bits_xcpt_ae_inst ; 
    wire core_ibuf_xcpt_1_pf_inst = core_ibuf_bufMask [1] ?  core_ibuf_buf_xcpt_pf_inst : core_ibuf_io_imem_bits_xcpt_pf_inst ; 
    wire core_ibuf_xcpt_1_gf_inst = core_ibuf_bufMask [1] ?  core_ibuf_buf_xcpt_gf_inst : core_ibuf_io_imem_bits_xcpt_gf_inst ; 
    wire core_ibuf_xcpt_1_ae_inst = core_ibuf_bufMask [1] ?  core_ibuf_buf_xcpt_ae_inst : core_ibuf_io_imem_bits_xcpt_ae_inst ; 
    wire[1:0] core_ibuf_buf_replay_0 = core_ibuf_buf_replay  ?  core_ibuf_bufMask :2'h0; 
    wire[1:0] core_ibuf_ic_replay = core_ibuf_buf_replay_0 |( core_ibuf_io_imem_bits_replay  ?  core_ibuf_valid &~ core_ibuf_bufMask :2'h0); 
  always @( posedge  core_ibuf_clock )
         begin 
             if (~ core_ibuf_reset &~(~ core_ibuf_io_imem_valid |~ core_ibuf_io_imem_bits_btb_taken | core_ibuf_io_imem_bits_btb_bridx >= core_ibuf_pcWordBits ))
                 begin 
                     if (1)$error("Assertion failed\n    at IBuf.scala:79 assert(!io.imem.valid || !io.imem.bits.btb.taken || io.imem.bits.btb.bridx >= pcWordBits)\n");
                     if (1)$fatal;
                 end 
         end
    wire core_ibuf_replay = core_ibuf_ic_replay [0]|~ core_ibuf__exp_io_rvc & core_ibuf_ic_replay [1]; 
    wire core_ibuf_full_insn = core_ibuf__exp_io_rvc | core_ibuf_valid [1]| core_ibuf_buf_replay_0 [0]; 
    wire[1:0] core_ibuf_io_inst_0_bits_xcpt1_hi ={ core_ibuf_xcpt_1_pf_inst , core_ibuf_xcpt_1_gf_inst }; 
    wire[2:0] core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 = core_ibuf__exp_io_rvc  ? 3'h0:{ core_ibuf_io_inst_0_bits_xcpt1_hi , core_ibuf_xcpt_1_ae_inst }; 
    wire core_ibuf__GEN_1 = core_ibuf_bufMask [0]& core_ibuf__exp_io_rvc | core_ibuf_bufMask [1]; 
  assign  core_ibuf_nReady = core_ibuf_full_insn  ? ( core_ibuf__exp_io_rvc  ? 2'h1:2'h2):2'h0; 
    wire[63:0] core_ibuf__buf_data_T_1 = core_ibuf_buf_data_data >>{58'h0, core_ibuf_shamt ,4'h0}; 
    wire core_ibuf__GEN_2 = core_ibuf_io_imem_valid & core_ibuf__nBufValid_T & core_ibuf_nICReady < core_ibuf_nIC &~( core_ibuf__nBufValid_T_6 [1]); 
  always @( posedge  core_ibuf_clock )
         begin 
             if ( core_ibuf_reset ) 
                 core_ibuf_nBufValid  <=1'h0;
              else  
                 core_ibuf_nBufValid  <=~ core_ibuf_io_kill &( core_ibuf_io_inst_0_ready  ? ( core_ibuf__GEN_2  ?  core_ibuf__nBufValid_T_6 [0]:~( core_ibuf__nBufValid_T |~ core_ibuf_nBufValid )& core_ibuf_nBufValid - core_ibuf_nReady [0]): core_ibuf_nBufValid );
             if ( core_ibuf_io_inst_0_ready & core_ibuf__GEN_2 )
                 begin  
                     core_ibuf_buf_btb_cfiType  <= core_ibuf_io_imem_bits_btb_cfiType ; 
                     core_ibuf_buf_btb_taken  <= core_ibuf_io_imem_bits_btb_taken ; 
                     core_ibuf_buf_btb_mask  <= core_ibuf_io_imem_bits_btb_mask ; 
                     core_ibuf_buf_btb_bridx  <= core_ibuf_io_imem_bits_btb_bridx ; 
                     core_ibuf_buf_btb_target  <= core_ibuf_io_imem_bits_btb_target ; 
                     core_ibuf_buf_btb_entry  <= core_ibuf_io_imem_bits_btb_entry ; 
                     core_ibuf_buf_btb_bht_history  <= core_ibuf_io_imem_bits_btb_bht_history ; 
                     core_ibuf_buf_btb_bht_value  <= core_ibuf_io_imem_bits_btb_bht_value ; 
                     core_ibuf_buf_pc  <= core_ibuf_io_imem_bits_pc &32'hFFFFFFFC| core_ibuf_io_imem_bits_pc +{29'h0, core_ibuf_nICReady ,1'h0}&32'h3; 
                     core_ibuf_buf_data  <={16'h0, core_ibuf__buf_data_T_1 [15:0]}; 
                     core_ibuf_buf_mask  <= core_ibuf_io_imem_bits_mask ; 
                     core_ibuf_buf_xcpt_pf_inst  <= core_ibuf_io_imem_bits_xcpt_pf_inst ; 
                     core_ibuf_buf_xcpt_gf_inst  <= core_ibuf_io_imem_bits_xcpt_gf_inst ; 
                     core_ibuf_buf_xcpt_ae_inst  <= core_ibuf_io_imem_bits_xcpt_ae_inst ; 
                     core_ibuf_buf_replay  <= core_ibuf_io_imem_bits_replay ; 
                     core_ibuf_ibufBTBResp_cfiType  <= core_ibuf_io_imem_bits_btb_cfiType ; 
                     core_ibuf_ibufBTBResp_taken  <= core_ibuf_io_imem_bits_btb_taken ; 
                     core_ibuf_ibufBTBResp_mask  <= core_ibuf_io_imem_bits_btb_mask ; 
                     core_ibuf_ibufBTBResp_bridx  <= core_ibuf_io_imem_bits_btb_bridx ; 
                     core_ibuf_ibufBTBResp_target  <= core_ibuf_io_imem_bits_btb_target ; 
                     core_ibuf_ibufBTBResp_entry  <= core_ibuf_io_imem_bits_btb_entry ; 
                     core_ibuf_ibufBTBResp_bht_history  <= core_ibuf_io_imem_bits_btb_bht_history ; 
                     core_ibuf_ibufBTBResp_bht_value  <= core_ibuf_io_imem_bits_btb_bht_value ;
                 end 
         end
    wire[31:0] core_ibuf_exp_io_in;
    wire[31:0] core_ibuf_exp_io_out_bits;
    wire[4:0] core_ibuf_exp_io_out_rd;
    wire[4:0] core_ibuf_exp_io_out_rs1;
    wire[4:0] core_ibuf_exp_io_out_rs2;
    wire[4:0] core_ibuf_exp_io_out_rs3;
    wire core_ibuf_exp_io_rvc;

    wire[31:0] core_ibuf_exp_io_out_s_24_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_25_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_26_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_27_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_28_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_29_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_30_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_31_bits = core_ibuf_exp_io_in ; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rd =5'h1; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rd =5'h1; 
    wire[11:0] core_ibuf_exp_io_out_s_jr_lo =12'h67; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rs1 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rd =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rs2 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rd =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rs2 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rs1 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rd =5'h0; 
    wire[11:0] core_ibuf_exp_io_out_s_jalr_lo =12'hE7; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rs1 =5'h2; 
    wire[6:0] core_ibuf_exp_io_out_s_opc =(|( core_ibuf_exp_io_in [12:5])) ? 7'h13:7'h1F; 
    wire[2:0] core_ibuf_exp__GEN ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[2:0] core_ibuf_exp_io_out_s_lo ; 
  assign  core_ibuf_exp_io_out_s_lo = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_3 ; 
  assign  core_ibuf_exp_io_out_s_lo_3 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_5 ; 
  assign  core_ibuf_exp_io_out_s_lo_5 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_7 ; 
  assign  core_ibuf_exp_io_out_s_lo_7 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_8 ; 
  assign  core_ibuf_exp_io_out_s_lo_8 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_11 ; 
  assign  core_ibuf_exp_io_out_s_lo_11 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_12 ; 
  assign  core_ibuf_exp_io_out_s_lo_12 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_14 ; 
  assign  core_ibuf_exp_io_out_s_lo_14 = core_ibuf_exp__GEN ; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_15 ; 
  assign  core_ibuf_exp_io_out_s_lo_15 = core_ibuf_exp__GEN ; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_hi ={ core_ibuf_exp_io_in [10:7], core_ibuf_exp_io_in [12:11]}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi ={ core_ibuf_exp_io_out_s_hi_hi , core_ibuf_exp_io_in [5]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_1 ={2'h1, core_ibuf_exp_io_in [4:2], core_ibuf_exp_io_out_s_opc }; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_hi_1 ={ core_ibuf_exp_io_out_s_hi , core_ibuf_exp_io_out_s_lo ,5'h2}; 
    wire[17:0] core_ibuf_exp_io_out_s_hi_1 ={ core_ibuf_exp_io_out_s_hi_hi_1 ,3'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_0_bits ={2'h0, core_ibuf_exp_io_out_s_hi_1 , core_ibuf_exp_io_out_s_lo_1 }; 
    wire[4:0] core_ibuf_exp__GEN_0 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_2 ; 
  assign  core_ibuf_exp_io_out_s_hi_2 = core_ibuf_exp__GEN_0 ; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_11 ; 
  assign  core_ibuf_exp_io_out_s_hi_11 = core_ibuf_exp__GEN_0 ; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_12 ; 
  assign  core_ibuf_exp_io_out_s_hi_12 = core_ibuf_exp__GEN_0 ; 
    wire[11:0] core_ibuf_exp__GEN_1 ={2'h1, core_ibuf_exp_io_in [4:2],7'h7}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_2 ; 
  assign  core_ibuf_exp_io_out_s_lo_2 = core_ibuf_exp__GEN_1 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_6 ; 
  assign  core_ibuf_exp_io_out_s_lo_6 = core_ibuf_exp__GEN_1 ; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_2 ={ core_ibuf_exp_io_out_s_hi_2 ,5'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[15:0] core_ibuf_exp_io_out_s_hi_3 ={ core_ibuf_exp_io_out_s_hi_hi_2 ,3'h3}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_1_bits ={4'h0, core_ibuf_exp_io_out_s_hi_3 , core_ibuf_exp_io_out_s_lo_2 }; 
    wire[3:0] core_ibuf_exp__GEN_2 ={ core_ibuf_exp_io_in [5], core_ibuf_exp_io_in [12:10]}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_4 ; 
  assign  core_ibuf_exp_io_out_s_hi_4 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_6 ; 
  assign  core_ibuf_exp_io_out_s_hi_6 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_8 ; 
  assign  core_ibuf_exp_io_out_s_hi_8 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_9 ; 
  assign  core_ibuf_exp_io_out_s_hi_9 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_14 ; 
  assign  core_ibuf_exp_io_out_s_hi_14 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_15 ; 
  assign  core_ibuf_exp_io_out_s_hi_15 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_17 ; 
  assign  core_ibuf_exp_io_out_s_hi_17 = core_ibuf_exp__GEN_2 ; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_18 ; 
  assign  core_ibuf_exp_io_out_s_hi_18 = core_ibuf_exp__GEN_2 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_4 ={2'h1, core_ibuf_exp_io_in [4:2],7'h3}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_hi_3 ={ core_ibuf_exp_io_out_s_hi_4 , core_ibuf_exp_io_out_s_lo_3 ,2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_5 ={ core_ibuf_exp_io_out_s_hi_hi_3 ,3'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_2_bits ={5'h0, core_ibuf_exp_io_out_s_hi_5 , core_ibuf_exp_io_out_s_lo_4 }; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_hi_4 ={ core_ibuf_exp_io_out_s_hi_6 , core_ibuf_exp_io_out_s_lo_5 ,2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_7 ={ core_ibuf_exp_io_out_s_hi_hi_4 ,3'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_3_bits ={5'h0, core_ibuf_exp_io_out_s_hi_7 , core_ibuf_exp_io_out_s_lo_6 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi ={3'h2, core_ibuf_exp_io_out_s_hi_9 [1:0], core_ibuf_exp_io_out_s_lo_8 }; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_9 ={ core_ibuf_exp_io_out_s_lo_hi ,7'h3F}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_5 ={ core_ibuf_exp_io_out_s_hi_8 [3:2],2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_10 ={ core_ibuf_exp_io_out_s_hi_hi_5 ,2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_4_bits ={5'h0, core_ibuf_exp_io_out_s_hi_10 , core_ibuf_exp_io_out_s_lo_9 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_1 ={3'h3, core_ibuf_exp_io_out_s_hi_12 [1:0],3'h0}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_10 ={ core_ibuf_exp_io_out_s_lo_hi_1 ,7'h27}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_hi_6 ={ core_ibuf_exp_io_out_s_hi_11 [4:2],2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_13 ={ core_ibuf_exp_io_out_s_hi_hi_6 ,2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_5_bits ={4'h0, core_ibuf_exp_io_out_s_hi_13 , core_ibuf_exp_io_out_s_lo_10 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_2 ={3'h2, core_ibuf_exp_io_out_s_hi_15 [1:0], core_ibuf_exp_io_out_s_lo_12 }; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_13 ={ core_ibuf_exp_io_out_s_lo_hi_2 ,7'h23}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_7 ={ core_ibuf_exp_io_out_s_hi_14 [3:2],2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_16 ={ core_ibuf_exp_io_out_s_hi_hi_7 ,2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_6_bits ={5'h0, core_ibuf_exp_io_out_s_hi_16 , core_ibuf_exp_io_out_s_lo_13 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_3 ={3'h2, core_ibuf_exp_io_out_s_hi_18 [1:0], core_ibuf_exp_io_out_s_lo_15 }; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_16 ={ core_ibuf_exp_io_out_s_lo_hi_3 ,7'h27}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_8 ={ core_ibuf_exp_io_out_s_hi_17 [3:2],2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_19 ={ core_ibuf_exp_io_out_s_hi_hi_8 ,2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_7_bits ={5'h0, core_ibuf_exp_io_out_s_hi_19 , core_ibuf_exp_io_out_s_lo_16 }; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rd = core_ibuf_exp_io_in [11:7]; 
    wire[11:0] core_ibuf_exp__GEN_3 ={ core_ibuf_exp_io_in [11:7],7'h13}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_17 ; 
  assign  core_ibuf_exp_io_out_s_lo_17 = core_ibuf_exp__GEN_3 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_23 ; 
  assign  core_ibuf_exp_io_out_s_lo_23 = core_ibuf_exp__GEN_3 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_45 ; 
  assign  core_ibuf_exp_io_out_s_lo_45 = core_ibuf_exp__GEN_3 ; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_9 ={{7{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:2], core_ibuf_exp_io_in [11:7]}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_20 ={ core_ibuf_exp_io_out_s_hi_hi_9 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_8_bits ={ core_ibuf_exp_io_out_s_hi_20 , core_ibuf_exp_io_out_s_lo_17 }; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[3:0] core_ibuf_exp__GEN_4 ={ core_ibuf_exp_io_in [5:3],1'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo ; 
  assign  core_ibuf_exp_io_out_s_lo_lo = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_1 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_1 = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_2 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_2 = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_3 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_3 = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_4 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_4 = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_5 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_5 = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_6 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_6 = core_ibuf_exp__GEN_4 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_7 ; 
  assign  core_ibuf_exp_io_out_s_lo_lo_7 = core_ibuf_exp__GEN_4 ; 
    wire[1:0] core_ibuf_exp__GEN_5 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [11]}; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_4 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_4 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_5 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_5 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_6 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_6 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_7 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_7 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_10 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_10 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_11 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_11 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_12 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_12 = core_ibuf_exp__GEN_5 ; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_13 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_13 = core_ibuf_exp__GEN_5 ; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_18 ={ core_ibuf_exp_io_out_s_lo_hi_4 , core_ibuf_exp_io_out_s_lo_lo }; 
    wire[1:0] core_ibuf_exp__GEN_6 ={ core_ibuf_exp_io_in [6], core_ibuf_exp_io_in [7]}; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo ; 
  assign  core_ibuf_exp_io_out_s_hi_lo = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_1 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_1 = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_2 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_2 = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_3 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_3 = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_4 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_4 = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_5 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_5 = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_6 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_6 = core_ibuf_exp__GEN_6 ; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_7 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_7 = core_ibuf_exp__GEN_6 ; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_10 ={ core_ibuf_exp_io_out_s_hi_hi_hi , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_21 ={ core_ibuf_exp_io_out_s_hi_hi_10 , core_ibuf_exp_io_out_s_hi_lo }; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_19 ={ core_ibuf_exp_io_out_s_lo_hi_5 , core_ibuf_exp_io_out_s_lo_lo_1 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_1 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_11 ={ core_ibuf_exp_io_out_s_hi_hi_hi_1 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_22 ={ core_ibuf_exp_io_out_s_hi_hi_11 , core_ibuf_exp_io_out_s_hi_lo_1 }; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_20 ={ core_ibuf_exp_io_out_s_lo_hi_6 , core_ibuf_exp_io_out_s_lo_lo_2 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_2 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_12 ={ core_ibuf_exp_io_out_s_hi_hi_hi_2 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_23 ={ core_ibuf_exp_io_out_s_hi_hi_12 , core_ibuf_exp_io_out_s_hi_lo_2 }; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_21 ={ core_ibuf_exp_io_out_s_lo_hi_7 , core_ibuf_exp_io_out_s_lo_lo_3 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_3 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_13 ={ core_ibuf_exp_io_out_s_hi_hi_hi_3 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_24 ={ core_ibuf_exp_io_out_s_hi_hi_13 , core_ibuf_exp_io_out_s_hi_lo_3 }; 
    wire[12:0] core_ibuf_exp_io_out_s_lo_hi_8 ={ core_ibuf_exp_io_out_s_hi_24 [13:6],5'h1}; 
    wire[19:0] core_ibuf_exp_io_out_s_lo_22 ={ core_ibuf_exp_io_out_s_lo_hi_8 ,7'h6F}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_14 ={ core_ibuf_exp_io_out_s_hi_21 [14], core_ibuf_exp_io_out_s_hi_22 [4:0], core_ibuf_exp_io_out_s_lo_19 [5:1]}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_25 ={ core_ibuf_exp_io_out_s_hi_hi_14 , core_ibuf_exp_io_out_s_hi_23 [5]}; 
    wire[31:0] core_ibuf_exp_io_out_s_9_bits ={ core_ibuf_exp_io_out_s_hi_25 , core_ibuf_exp_io_out_s_lo_22 }; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_15 ={{7{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:2],5'h0}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_26 ={ core_ibuf_exp_io_out_s_hi_hi_15 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_10_bits ={ core_ibuf_exp_io_out_s_hi_26 , core_ibuf_exp_io_out_s_lo_23 }; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_1 ={3'h3,{{7{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:2]}==12'h0,3'h7}; 
    wire[19:0] core_ibuf_exp_io_out_s_me_hi ={{15{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:2]}; 
    wire[24:0] core_ibuf_exp_io_out_s_me_hi_1 ={ core_ibuf_exp_io_out_s_me_hi , core_ibuf_exp_io_in [11:7]}; 
    wire[31:0] core_ibuf_exp_io_out_s_me_bits ={ core_ibuf_exp_io_out_s_me_hi_1 , core_ibuf_exp_io_out_s_opc_1 }; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire core_ibuf_exp__io_out_s_T_227 = core_ibuf_exp_io_in [11:7]==5'h0| core_ibuf_exp_io_in [11:7]==5'h2; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_2 =(|{{7{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:2]}) ? 7'h13:7'h1F; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_9 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [6]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_24 ={ core_ibuf_exp_io_out_s_lo_hi_9 ,4'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_hi_16 ={{3{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [4:3]}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_27 ={ core_ibuf_exp_io_out_s_hi_hi_16 , core_ibuf_exp_io_in [5]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_25 ={ core_ibuf_exp_io_in [11:7], core_ibuf_exp_io_out_s_opc_2 }; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_17 ={ core_ibuf_exp_io_out_s_hi_27 , core_ibuf_exp_io_out_s_lo_24 , core_ibuf_exp_io_in [11:7]}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_28 ={ core_ibuf_exp_io_out_s_hi_hi_17 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_res_bits ={ core_ibuf_exp_io_out_s_hi_28 , core_ibuf_exp_io_out_s_lo_25 }; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[31:0] core_ibuf_exp_io_out_s_11_bits = core_ibuf_exp__io_out_s_T_227  ?  core_ibuf_exp_io_out_s_res_bits : core_ibuf_exp_io_out_s_me_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rd = core_ibuf_exp__io_out_s_T_227  ?  core_ibuf_exp_io_out_s_res_rd : core_ibuf_exp_io_out_s_me_rd ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rs1 = core_ibuf_exp__io_out_s_T_227  ?  core_ibuf_exp_io_out_s_res_rs1 : core_ibuf_exp_io_out_s_me_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rs2 = core_ibuf_exp__io_out_s_T_227  ?  core_ibuf_exp_io_out_s_res_rs2 : core_ibuf_exp_io_out_s_me_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rs3 = core_ibuf_exp__io_out_s_T_227  ?  core_ibuf_exp_io_out_s_res_rs3 : core_ibuf_exp_io_out_s_me_rs3 ; 
    wire[11:0] core_ibuf_exp__GEN_7 ={2'h1, core_ibuf_exp_io_in [9:7],7'h13}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_26 ; 
  assign  core_ibuf_exp_io_out_s_lo_26 = core_ibuf_exp__GEN_7 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_27 ; 
  assign  core_ibuf_exp_io_out_s_lo_27 = core_ibuf_exp__GEN_7 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_28 ; 
  assign  core_ibuf_exp_io_out_s_lo_28 = core_ibuf_exp__GEN_7 ; 
    wire[10:0] core_ibuf_exp__GEN_8 ={ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:2],2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_18 ; 
  assign  core_ibuf_exp_io_out_s_hi_hi_18 = core_ibuf_exp__GEN_8 ; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_19 ; 
  assign  core_ibuf_exp_io_out_s_hi_hi_19 = core_ibuf_exp__GEN_8 ; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_29 ={ core_ibuf_exp_io_out_s_hi_hi_18 ,3'h5}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_30 ={ core_ibuf_exp_io_out_s_hi_hi_19 ,3'h5}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_20 ={{7{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:2],2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_31 ={ core_ibuf_exp_io_out_s_hi_hi_20 ,3'h7}; reg[2:0] core_ibuf_exp_casez_tmp ; 
    wire[2:0] core_ibuf_exp__io_out_s_funct_T_2 ={ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:5]}; 
    wire[2:0] core_ibuf_exp__io_out_s_funct_T_4 ={ core_ibuf_exp__io_out_s_funct_T_2 ==3'h1,2'h0}; 
  always @(*)
         begin 
             casez ( core_ibuf_exp__io_out_s_funct_T_2 )
              3 'b000: 
                  core_ibuf_exp_casez_tmp  = core_ibuf_exp__io_out_s_funct_T_4 ;
              3 'b001: 
                  core_ibuf_exp_casez_tmp  = core_ibuf_exp__io_out_s_funct_T_4 ;
              3 'b010: 
                  core_ibuf_exp_casez_tmp  =3'h6;
              3 'b011: 
                  core_ibuf_exp_casez_tmp  =3'h7;
              3 'b100: 
                  core_ibuf_exp_casez_tmp  =3'h0;
              3 'b101: 
                  core_ibuf_exp_casez_tmp  =3'h0;
              3 'b110: 
                  core_ibuf_exp_casez_tmp  =3'h2;
              default : 
                  core_ibuf_exp_casez_tmp  =3'h3;endcase
         end
    wire[2:0] core_ibuf_exp_io_out_s_funct = core_ibuf_exp_casez_tmp ; 
    wire[30:0] core_ibuf_exp_io_out_s_sub ={ core_ibuf_exp_io_in [6:5]==2'h0,30'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_3 ={3'h3, core_ibuf_exp_io_in [12],3'h3}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_29 ={2'h1, core_ibuf_exp_io_in [9:7], core_ibuf_exp_io_out_s_opc_3 }; 
    wire[9:0] core_ibuf_exp_io_out_s_hi_hi_21 ={2'h1, core_ibuf_exp_io_in [4:2],2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_32 ={ core_ibuf_exp_io_out_s_hi_hi_21 , core_ibuf_exp_io_out_s_funct }; 
    wire[31:0] core_ibuf_exp_io_out_s_12_bits =(&( core_ibuf_exp_io_in [11:10])) ? {1'h0,{6'h0, core_ibuf_exp_io_out_s_hi_32 , core_ibuf_exp_io_out_s_lo_29 }| core_ibuf_exp_io_out_s_sub }: core_ibuf_exp_io_in [11:10]==2'h2 ? { core_ibuf_exp_io_out_s_hi_31 , core_ibuf_exp_io_out_s_lo_28 }:{1'h0, core_ibuf_exp_io_in [11:10]==2'h1 ? {5'h10, core_ibuf_exp_io_out_s_hi_30 , core_ibuf_exp_io_out_s_lo_27 }:{5'h0, core_ibuf_exp_io_out_s_hi_29 , core_ibuf_exp_io_out_s_lo_26 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rd ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_30 ={ core_ibuf_exp_io_out_s_lo_hi_10 , core_ibuf_exp_io_out_s_lo_lo_4 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_4 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_22 ={ core_ibuf_exp_io_out_s_hi_hi_hi_4 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_33 ={ core_ibuf_exp_io_out_s_hi_hi_22 , core_ibuf_exp_io_out_s_hi_lo_4 }; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_31 ={ core_ibuf_exp_io_out_s_lo_hi_11 , core_ibuf_exp_io_out_s_lo_lo_5 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_5 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_23 ={ core_ibuf_exp_io_out_s_hi_hi_hi_5 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_34 ={ core_ibuf_exp_io_out_s_hi_hi_23 , core_ibuf_exp_io_out_s_hi_lo_5 }; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_32 ={ core_ibuf_exp_io_out_s_lo_hi_12 , core_ibuf_exp_io_out_s_lo_lo_6 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_6 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_24 ={ core_ibuf_exp_io_out_s_hi_hi_hi_6 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_35 ={ core_ibuf_exp_io_out_s_hi_hi_24 , core_ibuf_exp_io_out_s_hi_lo_6 }; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_33 ={ core_ibuf_exp_io_out_s_lo_hi_13 , core_ibuf_exp_io_out_s_lo_lo_7 }; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_7 ={{10{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_25 ={ core_ibuf_exp_io_out_s_hi_hi_hi_7 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_36 ={ core_ibuf_exp_io_out_s_hi_hi_25 , core_ibuf_exp_io_out_s_hi_lo_7 }; 
    wire[12:0] core_ibuf_exp_io_out_s_lo_hi_14 ={ core_ibuf_exp_io_out_s_hi_36 [13:6],5'h0}; 
    wire[19:0] core_ibuf_exp_io_out_s_lo_34 ={ core_ibuf_exp_io_out_s_lo_hi_14 ,7'h6F}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_26 ={ core_ibuf_exp_io_out_s_hi_33 [14], core_ibuf_exp_io_out_s_hi_34 [4:0], core_ibuf_exp_io_out_s_lo_31 [5:1]}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_37 ={ core_ibuf_exp_io_out_s_hi_hi_26 , core_ibuf_exp_io_out_s_hi_35 [5]}; 
    wire[31:0] core_ibuf_exp_io_out_s_13_bits ={ core_ibuf_exp_io_out_s_hi_37 , core_ibuf_exp_io_out_s_lo_34 }; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[3:0] core_ibuf_exp__GEN_9 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_15 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_15 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_16 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_16 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_17 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_17 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_18 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_18 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_20 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_20 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_21 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_21 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_22 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_22 = core_ibuf_exp__GEN_9 ; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_23 ; 
  assign  core_ibuf_exp_io_out_s_lo_hi_23 = core_ibuf_exp__GEN_9 ; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_35 ={ core_ibuf_exp_io_out_s_lo_hi_15 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_27 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_38 ={ core_ibuf_exp_io_out_s_hi_hi_27 , core_ibuf_exp_io_in [2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_36 ={ core_ibuf_exp_io_out_s_lo_hi_16 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_28 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_39 ={ core_ibuf_exp_io_out_s_hi_hi_28 , core_ibuf_exp_io_in [2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_37 ={ core_ibuf_exp_io_out_s_lo_hi_17 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_29 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_40 ={ core_ibuf_exp_io_out_s_hi_hi_29 , core_ibuf_exp_io_in [2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_38 ={ core_ibuf_exp_io_out_s_lo_hi_18 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_30 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_41 ={ core_ibuf_exp_io_out_s_hi_hi_30 , core_ibuf_exp_io_in [2]}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_lo_8 ={ core_ibuf_exp_io_out_s_hi_41 [6],7'h63}; 
    wire[6:0] core_ibuf_exp_io_out_s_lo_hi_19 ={3'h0, core_ibuf_exp_io_out_s_lo_37 [4:1]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_39 ={ core_ibuf_exp_io_out_s_lo_hi_19 , core_ibuf_exp_io_out_s_lo_lo_8 }; 
    wire[9:0] core_ibuf_exp__GEN_10 ={7'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[9:0] core_ibuf_exp_io_out_s_hi_lo_8 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_8 = core_ibuf_exp__GEN_10 ; 
    wire[9:0] core_ibuf_exp_io_out_s_hi_lo_9 ; 
  assign  core_ibuf_exp_io_out_s_hi_lo_9 = core_ibuf_exp__GEN_10 ; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_31 ={ core_ibuf_exp_io_out_s_hi_38 [7], core_ibuf_exp_io_out_s_hi_39 [5:0]}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_42 ={ core_ibuf_exp_io_out_s_hi_hi_31 , core_ibuf_exp_io_out_s_hi_lo_8 }; 
    wire[31:0] core_ibuf_exp_io_out_s_14_bits ={ core_ibuf_exp_io_out_s_hi_42 , core_ibuf_exp_io_out_s_lo_39 }; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rd ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_40 ={ core_ibuf_exp_io_out_s_lo_hi_20 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_32 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_43 ={ core_ibuf_exp_io_out_s_hi_hi_32 , core_ibuf_exp_io_in [2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_41 ={ core_ibuf_exp_io_out_s_lo_hi_21 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_33 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_44 ={ core_ibuf_exp_io_out_s_hi_hi_33 , core_ibuf_exp_io_in [2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_42 ={ core_ibuf_exp_io_out_s_lo_hi_22 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_34 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_45 ={ core_ibuf_exp_io_out_s_hi_hi_34 , core_ibuf_exp_io_in [2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_43 ={ core_ibuf_exp_io_out_s_lo_hi_23 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_35 ={{5{ core_ibuf_exp_io_in [12]}}, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_46 ={ core_ibuf_exp_io_out_s_hi_hi_35 , core_ibuf_exp_io_in [2]}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_lo_9 ={ core_ibuf_exp_io_out_s_hi_46 [6],7'h63}; 
    wire[6:0] core_ibuf_exp_io_out_s_lo_hi_24 ={3'h1, core_ibuf_exp_io_out_s_lo_42 [4:1]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_44 ={ core_ibuf_exp_io_out_s_lo_hi_24 , core_ibuf_exp_io_out_s_lo_lo_9 }; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_36 ={ core_ibuf_exp_io_out_s_hi_43 [7], core_ibuf_exp_io_out_s_hi_44 [5:0]}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_47 ={ core_ibuf_exp_io_out_s_hi_hi_36 , core_ibuf_exp_io_out_s_hi_lo_9 }; 
    wire[31:0] core_ibuf_exp_io_out_s_15_bits ={ core_ibuf_exp_io_out_s_hi_47 , core_ibuf_exp_io_out_s_lo_44 }; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[6:0] core_ibuf_exp_io_out_s_load_opc =(|( core_ibuf_exp_io_in [11:7])) ? 7'h3:7'h1F; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_37 ={ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:2], core_ibuf_exp_io_in [11:7]}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_48 ={ core_ibuf_exp_io_out_s_hi_hi_37 ,3'h1}; 
    wire[31:0] core_ibuf_exp_io_out_s_16_bits ={6'h0, core_ibuf_exp_io_out_s_hi_48 , core_ibuf_exp_io_out_s_lo_45 }; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_46 ={ core_ibuf_exp_io_in [6:5],3'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_49 ={ core_ibuf_exp_io_in [4:2], core_ibuf_exp_io_in [12]}; 
    wire[11:0] core_ibuf_exp__GEN_11 ={ core_ibuf_exp_io_in [11:7],7'h7}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_47 ; 
  assign  core_ibuf_exp_io_out_s_lo_47 = core_ibuf_exp__GEN_11 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_51 ; 
  assign  core_ibuf_exp_io_out_s_lo_51 = core_ibuf_exp__GEN_11 ; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_hi_38 ={ core_ibuf_exp_io_out_s_hi_49 , core_ibuf_exp_io_out_s_lo_46 ,5'h2}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_50 ={ core_ibuf_exp_io_out_s_hi_hi_38 ,3'h3}; 
    wire[31:0] core_ibuf_exp_io_out_s_17_bits ={3'h0, core_ibuf_exp_io_out_s_hi_50 , core_ibuf_exp_io_out_s_lo_47 }; 
    wire[4:0] core_ibuf_exp__GEN_12 ={ core_ibuf_exp_io_in [6:4],2'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_48 ; 
  assign  core_ibuf_exp_io_out_s_lo_48 = core_ibuf_exp__GEN_12 ; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_50 ; 
  assign  core_ibuf_exp_io_out_s_lo_50 = core_ibuf_exp__GEN_12 ; 
    wire[2:0] core_ibuf_exp__GEN_13 ={ core_ibuf_exp_io_in [3:2], core_ibuf_exp_io_in [12]}; 
    wire[2:0] core_ibuf_exp_io_out_s_hi_51 ; 
  assign  core_ibuf_exp_io_out_s_hi_51 = core_ibuf_exp__GEN_13 ; 
    wire[2:0] core_ibuf_exp_io_out_s_hi_53 ; 
  assign  core_ibuf_exp_io_out_s_hi_53 = core_ibuf_exp__GEN_13 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_49 ={ core_ibuf_exp_io_in [11:7], core_ibuf_exp_io_out_s_load_opc }; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_39 ={ core_ibuf_exp_io_out_s_hi_51 , core_ibuf_exp_io_out_s_lo_48 ,5'h2}; 
    wire[15:0] core_ibuf_exp_io_out_s_hi_52 ={ core_ibuf_exp_io_out_s_hi_hi_39 ,3'h2}; 
    wire[31:0] core_ibuf_exp_io_out_s_18_bits ={4'h0, core_ibuf_exp_io_out_s_hi_52 , core_ibuf_exp_io_out_s_lo_49 }; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_40 ={ core_ibuf_exp_io_out_s_hi_53 , core_ibuf_exp_io_out_s_lo_50 ,5'h2}; 
    wire[15:0] core_ibuf_exp_io_out_s_hi_54 ={ core_ibuf_exp_io_out_s_hi_hi_40 ,3'h2}; 
    wire[31:0] core_ibuf_exp_io_out_s_19_bits ={4'h0, core_ibuf_exp_io_out_s_hi_54 , core_ibuf_exp_io_out_s_lo_51 }; 
    wire[11:0] core_ibuf_exp__GEN_14 ={ core_ibuf_exp_io_in [11:7],7'h33}; 
    wire[11:0] core_ibuf_exp_io_out_s_mv_lo ; 
  assign  core_ibuf_exp_io_out_s_mv_lo = core_ibuf_exp__GEN_14 ; 
    wire[11:0] core_ibuf_exp_io_out_s_add_lo ; 
  assign  core_ibuf_exp_io_out_s_add_lo = core_ibuf_exp__GEN_14 ; 
    wire[9:0] core_ibuf_exp_io_out_s_mv_hi_hi ={ core_ibuf_exp_io_in [6:2],5'h0}; 
    wire[12:0] core_ibuf_exp_io_out_s_mv_hi ={ core_ibuf_exp_io_out_s_mv_hi_hi ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_mv_bits ={7'h0, core_ibuf_exp_io_out_s_mv_hi , core_ibuf_exp_io_out_s_mv_lo }; 
    wire[9:0] core_ibuf_exp__GEN_15 ={ core_ibuf_exp_io_in [6:2], core_ibuf_exp_io_in [11:7]}; 
    wire[9:0] core_ibuf_exp_io_out_s_add_hi_hi ; 
  assign  core_ibuf_exp_io_out_s_add_hi_hi = core_ibuf_exp__GEN_15 ; 
    wire[9:0] core_ibuf_exp_io_out_s_jr_hi_hi ; 
  assign  core_ibuf_exp_io_out_s_jr_hi_hi = core_ibuf_exp__GEN_15 ; 
    wire[9:0] core_ibuf_exp_io_out_s_jalr_hi_hi ; 
  assign  core_ibuf_exp_io_out_s_jalr_hi_hi = core_ibuf_exp__GEN_15 ; 
    wire[12:0] core_ibuf_exp_io_out_s_add_hi ={ core_ibuf_exp_io_out_s_add_hi_hi ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_add_bits ={7'h0, core_ibuf_exp_io_out_s_add_hi , core_ibuf_exp_io_out_s_add_lo }; 
    wire[12:0] core_ibuf_exp_io_out_s_jr_hi ={ core_ibuf_exp_io_out_s_jr_hi_hi ,3'h0}; 
    wire[24:0] core_ibuf_exp_io_out_s_jr ={ core_ibuf_exp_io_out_s_jr_hi ,12'h67}; 
    wire[24:0] core_ibuf_exp_io_out_s_reserved ={ core_ibuf_exp_io_out_s_jr [24:7],7'h1F}; 
    wire[31:0] core_ibuf_exp_io_out_s_jr_reserved_bits ={7'h0,(|( core_ibuf_exp_io_in [11:7])) ?  core_ibuf_exp_io_out_s_jr : core_ibuf_exp_io_out_s_reserved }; 
    wire[31:0] core_ibuf_exp_io_out_s_jr_mv_bits =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_mv_bits : core_ibuf_exp_io_out_s_jr_reserved_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rd =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_mv_rd :5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rs1 =(|( core_ibuf_exp_io_in [6:2])) ? 5'h0: core_ibuf_exp_io_out_s_jr_reserved_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rs2 =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_mv_rs2 : core_ibuf_exp_io_out_s_jr_reserved_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rs3 =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_mv_rs3 : core_ibuf_exp_io_out_s_jr_reserved_rs3 ; 
    wire[12:0] core_ibuf_exp_io_out_s_jalr_hi ={ core_ibuf_exp_io_out_s_jalr_hi_hi ,3'h0}; 
    wire[24:0] core_ibuf_exp_io_out_s_jalr ={ core_ibuf_exp_io_out_s_jalr_hi ,12'hE7}; 
    wire[24:0] core_ibuf_exp_io_out_s_ebreak ={ core_ibuf_exp_io_out_s_jr [24:21], core_ibuf_exp_io_out_s_jr [20:7]|14'h2000,7'h73}; 
    wire[31:0] core_ibuf_exp_io_out_s_jalr_ebreak_bits ={7'h0,(|( core_ibuf_exp_io_in [11:7])) ?  core_ibuf_exp_io_out_s_jalr : core_ibuf_exp_io_out_s_ebreak }; 
    wire[31:0] core_ibuf_exp_io_out_s_jalr_add_bits =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_add_bits : core_ibuf_exp_io_out_s_jalr_ebreak_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rd =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_add_rd :5'h1; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rs1 =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_add_rs1 : core_ibuf_exp_io_out_s_jalr_ebreak_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rs2 =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_add_rs2 : core_ibuf_exp_io_out_s_jalr_ebreak_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rs3 =(|( core_ibuf_exp_io_in [6:2])) ?  core_ibuf_exp_io_out_s_add_rs3 : core_ibuf_exp_io_out_s_jalr_ebreak_rs3 ; 
    wire[31:0] core_ibuf_exp_io_out_s_20_bits = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_bits : core_ibuf_exp_io_out_s_jr_mv_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rd = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rd : core_ibuf_exp_io_out_s_jr_mv_rd ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rs1 = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rs1 : core_ibuf_exp_io_out_s_jr_mv_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rs2 = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rs2 : core_ibuf_exp_io_out_s_jr_mv_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rs3 = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rs3 : core_ibuf_exp_io_out_s_jr_mv_rs3 ; 
    wire[5:0] core_ibuf_exp__GEN_16 ={ core_ibuf_exp_io_in [9:7], core_ibuf_exp_io_in [12:10]}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_55 ; 
  assign  core_ibuf_exp_io_out_s_hi_55 = core_ibuf_exp__GEN_16 ; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_56 ; 
  assign  core_ibuf_exp_io_out_s_hi_56 = core_ibuf_exp__GEN_16 ; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_25 ={3'h3, core_ibuf_exp_io_out_s_hi_56 [1:0],3'h0}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_52 ={ core_ibuf_exp_io_out_s_lo_hi_25 ,7'h27}; 
    wire[8:0] core_ibuf_exp_io_out_s_hi_hi_41 ={ core_ibuf_exp_io_out_s_hi_55 [5:2], core_ibuf_exp_io_in [6:2]}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_57 ={ core_ibuf_exp_io_out_s_hi_hi_41 ,5'h2}; 
    wire[31:0] core_ibuf_exp_io_out_s_21_bits ={3'h0, core_ibuf_exp_io_out_s_hi_57 , core_ibuf_exp_io_out_s_lo_52 }; 
    wire[5:0] core_ibuf_exp__GEN_17 ={ core_ibuf_exp_io_in [8:7], core_ibuf_exp_io_in [12:9]}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_58 ; 
  assign  core_ibuf_exp_io_out_s_hi_58 = core_ibuf_exp__GEN_17 ; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_59 ; 
  assign  core_ibuf_exp_io_out_s_hi_59 = core_ibuf_exp__GEN_17 ; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_61 ; 
  assign  core_ibuf_exp_io_out_s_hi_61 = core_ibuf_exp__GEN_17 ; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_62 ; 
  assign  core_ibuf_exp_io_out_s_hi_62 = core_ibuf_exp__GEN_17 ; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_26 ={3'h2, core_ibuf_exp_io_out_s_hi_59 [2:0],2'h0}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_53 ={ core_ibuf_exp_io_out_s_lo_hi_26 ,7'h23}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_hi_42 ={ core_ibuf_exp_io_out_s_hi_58 [5:3], core_ibuf_exp_io_in [6:2]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_60 ={ core_ibuf_exp_io_out_s_hi_hi_42 ,5'h2}; 
    wire[31:0] core_ibuf_exp_io_out_s_22_bits ={4'h0, core_ibuf_exp_io_out_s_hi_60 , core_ibuf_exp_io_out_s_lo_53 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_27 ={3'h2, core_ibuf_exp_io_out_s_hi_62 [2:0],2'h0}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_54 ={ core_ibuf_exp_io_out_s_lo_hi_27 ,7'h27}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_hi_43 ={ core_ibuf_exp_io_out_s_hi_61 [5:3], core_ibuf_exp_io_in [6:2]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_63 ={ core_ibuf_exp_io_out_s_hi_hi_43 ,5'h2}; 
    wire[31:0] core_ibuf_exp_io_out_s_23_bits ={4'h0, core_ibuf_exp_io_out_s_hi_63 , core_ibuf_exp_io_out_s_lo_54 }; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp__io_out_T_2 ={ core_ibuf_exp_io_in [1:0], core_ibuf_exp_io_in [15:13]}; reg[31:0] core_ibuf_exp_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( core_ibuf_exp__io_out_T_2 )
              5 'b00000: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_0_bits ;
              5 'b00001: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_1_bits ;
              5 'b00010: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_2_bits ;
              5 'b00011: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_3_bits ;
              5 'b00100: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_4_bits ;
              5 'b00101: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_5_bits ;
              5 'b00110: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_6_bits ;
              5 'b00111: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_7_bits ;
              5 'b01000: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_8_bits ;
              5 'b01001: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_9_bits ;
              5 'b01010: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_10_bits ;
              5 'b01011: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_11_bits ;
              5 'b01100: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_12_bits ;
              5 'b01101: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_13_bits ;
              5 'b01110: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_14_bits ;
              5 'b01111: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_15_bits ;
              5 'b10000: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_16_bits ;
              5 'b10001: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_17_bits ;
              5 'b10010: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_18_bits ;
              5 'b10011: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_19_bits ;
              5 'b10100: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_20_bits ;
              5 'b10101: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_21_bits ;
              5 'b10110: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_22_bits ;
              5 'b10111: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_23_bits ;
              5 'b11000: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_24_bits ;
              5 'b11001: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_25_bits ;
              5 'b11010: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_26_bits ;
              5 'b11011: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_27_bits ;
              5 'b11100: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_28_bits ;
              5 'b11101: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_29_bits ;
              5 'b11110: 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_30_bits ;
              default : 
                  core_ibuf_exp_casez_tmp_0  = core_ibuf_exp_io_out_s_31_bits ;endcase
         end
  reg[4:0] core_ibuf_exp_casez_tmp_1 ; 
  always @(*)
         begin 
             casez ( core_ibuf_exp__io_out_T_2 )
              5 'b00000: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_0_rd ;
              5 'b00001: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_1_rd ;
              5 'b00010: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_2_rd ;
              5 'b00011: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_3_rd ;
              5 'b00100: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_4_rd ;
              5 'b00101: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_5_rd ;
              5 'b00110: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_6_rd ;
              5 'b00111: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_7_rd ;
              5 'b01000: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_8_rd ;
              5 'b01001: 
                  core_ibuf_exp_casez_tmp_1  =5'h1;
              5 'b01010: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_10_rd ;
              5 'b01011: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_11_rd ;
              5 'b01100: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_12_rd ;
              5 'b01101: 
                  core_ibuf_exp_casez_tmp_1  =5'h0;
              5 'b01110: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_14_rd ;
              5 'b01111: 
                  core_ibuf_exp_casez_tmp_1  =5'h0;
              5 'b10000: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_16_rd ;
              5 'b10001: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_17_rd ;
              5 'b10010: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_18_rd ;
              5 'b10011: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_19_rd ;
              5 'b10100: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_20_rd ;
              5 'b10101: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_21_rd ;
              5 'b10110: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_22_rd ;
              5 'b10111: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_23_rd ;
              5 'b11000: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_24_rd ;
              5 'b11001: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_25_rd ;
              5 'b11010: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_26_rd ;
              5 'b11011: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_27_rd ;
              5 'b11100: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_28_rd ;
              5 'b11101: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_29_rd ;
              5 'b11110: 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_30_rd ;
              default : 
                  core_ibuf_exp_casez_tmp_1  = core_ibuf_exp_io_out_s_31_rd ;endcase
         end
  reg[4:0] core_ibuf_exp_casez_tmp_2 ; 
  always @(*)
         begin 
             casez ( core_ibuf_exp__io_out_T_2 )
              5 'b00000: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b00001: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_1_rs1 ;
              5 'b00010: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_2_rs1 ;
              5 'b00011: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_3_rs1 ;
              5 'b00100: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_4_rs1 ;
              5 'b00101: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_5_rs1 ;
              5 'b00110: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_6_rs1 ;
              5 'b00111: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_7_rs1 ;
              5 'b01000: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_8_rs1 ;
              5 'b01001: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_9_rs1 ;
              5 'b01010: 
                  core_ibuf_exp_casez_tmp_2  =5'h0;
              5 'b01011: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_11_rs1 ;
              5 'b01100: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_12_rs1 ;
              5 'b01101: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_13_rs1 ;
              5 'b01110: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_14_rs1 ;
              5 'b01111: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_15_rs1 ;
              5 'b10000: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_16_rs1 ;
              5 'b10001: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b10010: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b10011: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b10100: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_20_rs1 ;
              5 'b10101: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b10110: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b10111: 
                  core_ibuf_exp_casez_tmp_2  =5'h2;
              5 'b11000: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_24_rs1 ;
              5 'b11001: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_25_rs1 ;
              5 'b11010: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_26_rs1 ;
              5 'b11011: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_27_rs1 ;
              5 'b11100: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_28_rs1 ;
              5 'b11101: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_29_rs1 ;
              5 'b11110: 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_30_rs1 ;
              default : 
                  core_ibuf_exp_casez_tmp_2  = core_ibuf_exp_io_out_s_31_rs1 ;endcase
         end
  reg[4:0] core_ibuf_exp_casez_tmp_3 ; 
  always @(*)
         begin 
             casez ( core_ibuf_exp__io_out_T_2 )
              5 'b00000: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_0_rs2 ;
              5 'b00001: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_1_rs2 ;
              5 'b00010: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_2_rs2 ;
              5 'b00011: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_3_rs2 ;
              5 'b00100: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_4_rs2 ;
              5 'b00101: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_5_rs2 ;
              5 'b00110: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_6_rs2 ;
              5 'b00111: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_7_rs2 ;
              5 'b01000: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_8_rs2 ;
              5 'b01001: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_9_rs2 ;
              5 'b01010: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_10_rs2 ;
              5 'b01011: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_11_rs2 ;
              5 'b01100: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_12_rs2 ;
              5 'b01101: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_13_rs2 ;
              5 'b01110: 
                  core_ibuf_exp_casez_tmp_3  =5'h0;
              5 'b01111: 
                  core_ibuf_exp_casez_tmp_3  =5'h0;
              5 'b10000: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_16_rs2 ;
              5 'b10001: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_17_rs2 ;
              5 'b10010: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_18_rs2 ;
              5 'b10011: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_19_rs2 ;
              5 'b10100: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_20_rs2 ;
              5 'b10101: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_21_rs2 ;
              5 'b10110: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_22_rs2 ;
              5 'b10111: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_23_rs2 ;
              5 'b11000: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_24_rs2 ;
              5 'b11001: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_25_rs2 ;
              5 'b11010: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_26_rs2 ;
              5 'b11011: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_27_rs2 ;
              5 'b11100: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_28_rs2 ;
              5 'b11101: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_29_rs2 ;
              5 'b11110: 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_30_rs2 ;
              default : 
                  core_ibuf_exp_casez_tmp_3  = core_ibuf_exp_io_out_s_31_rs2 ;endcase
         end
  reg[4:0] core_ibuf_exp_casez_tmp_4 ; 
  always @(*)
         begin 
             casez ( core_ibuf_exp__io_out_T_2 )
              5 'b00000: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_0_rs3 ;
              5 'b00001: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_1_rs3 ;
              5 'b00010: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_2_rs3 ;
              5 'b00011: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_3_rs3 ;
              5 'b00100: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_4_rs3 ;
              5 'b00101: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_5_rs3 ;
              5 'b00110: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_6_rs3 ;
              5 'b00111: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_7_rs3 ;
              5 'b01000: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_8_rs3 ;
              5 'b01001: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_9_rs3 ;
              5 'b01010: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_10_rs3 ;
              5 'b01011: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_11_rs3 ;
              5 'b01100: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_12_rs3 ;
              5 'b01101: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_13_rs3 ;
              5 'b01110: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_14_rs3 ;
              5 'b01111: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_15_rs3 ;
              5 'b10000: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_16_rs3 ;
              5 'b10001: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_17_rs3 ;
              5 'b10010: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_18_rs3 ;
              5 'b10011: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_19_rs3 ;
              5 'b10100: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_20_rs3 ;
              5 'b10101: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_21_rs3 ;
              5 'b10110: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_22_rs3 ;
              5 'b10111: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_23_rs3 ;
              5 'b11000: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_24_rs3 ;
              5 'b11001: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_25_rs3 ;
              5 'b11010: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_26_rs3 ;
              5 'b11011: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_27_rs3 ;
              5 'b11100: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_28_rs3 ;
              5 'b11101: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_29_rs3 ;
              5 'b11110: 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_30_rs3 ;
              default : 
                  core_ibuf_exp_casez_tmp_4  = core_ibuf_exp_io_out_s_31_rs3 ;endcase
         end
  assign  core_ibuf_exp_io_out_bits = core_ibuf_exp_casez_tmp_0 ; 
  assign  core_ibuf_exp_io_out_rd = core_ibuf_exp_casez_tmp_1 ; 
  assign  core_ibuf_exp_io_out_rs1 = core_ibuf_exp_casez_tmp_2 ; 
  assign  core_ibuf_exp_io_out_rs2 = core_ibuf_exp_casez_tmp_3 ; 
  assign  core_ibuf_exp_io_out_rs3 = core_ibuf_exp_casez_tmp_4 ; 
  assign  core_ibuf_exp_io_rvc = core_ibuf_exp_io_in [1:0]!=2'h3;
    assign core_ibuf_exp_io_in = core_ibuf_inst;
    assign core_ibuf_io_inst_0_bits_inst_bits = core_ibuf_exp_io_out_bits;
    assign core_ibuf_io_inst_0_bits_inst_rd = core_ibuf_exp_io_out_rd;
    assign core_ibuf_io_inst_0_bits_inst_rs1 = core_ibuf_exp_io_out_rs1;
    assign core_ibuf_io_inst_0_bits_inst_rs2 = core_ibuf_exp_io_out_rs2;
    assign core_ibuf_io_inst_0_bits_inst_rs3 = core_ibuf_exp_io_out_rs3;
    assign core_ibuf__exp_io_rvc = core_ibuf_exp_io_rvc;
     
  assign  core_ibuf_io_imem_ready = core_ibuf_io_inst_0_ready & core_ibuf__nBufValid_T &( core_ibuf_nICReady >= core_ibuf_nIC |~( core_ibuf__nBufValid_T_6 [1])); 
  assign  core_ibuf_io_pc = core_ibuf_nBufValid  ?  core_ibuf_buf_pc : core_ibuf_io_imem_bits_pc ; 
  assign  core_ibuf_io_btb_resp_cfiType = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_cfiType : core_ibuf_io_imem_bits_btb_cfiType ; 
  assign  core_ibuf_io_btb_resp_taken = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_taken : core_ibuf_io_imem_bits_btb_taken ; 
  assign  core_ibuf_io_btb_resp_mask = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_mask : core_ibuf_io_imem_bits_btb_mask ; 
  assign  core_ibuf_io_btb_resp_bridx = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_bridx : core_ibuf_io_imem_bits_btb_bridx ; 
  assign  core_ibuf_io_btb_resp_target = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_target : core_ibuf_io_imem_bits_btb_target ; 
  assign  core_ibuf_io_btb_resp_entry = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_entry : core_ibuf_io_imem_bits_btb_entry ; 
  assign  core_ibuf_io_btb_resp_bht_history = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_bht_history : core_ibuf_io_imem_bits_btb_bht_history ; 
  assign  core_ibuf_io_btb_resp_bht_value = core_ibuf__GEN_1  ?  core_ibuf_ibufBTBResp_bht_value : core_ibuf_io_imem_bits_btb_bht_value ; 
  assign  core_ibuf_io_inst_0_valid = core_ibuf_valid [0]& core_ibuf_full_insn ; 
  assign  core_ibuf_io_inst_0_bits_xcpt0_pf_inst = core_ibuf_xcpt_0_pf_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt0_gf_inst = core_ibuf_xcpt_0_gf_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt0_ae_inst = core_ibuf_xcpt_0_ae_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt1_pf_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 [2]; 
  assign  core_ibuf_io_inst_0_bits_xcpt1_gf_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 [1]; 
  assign  core_ibuf_io_inst_0_bits_xcpt1_ae_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 [0]; 
  assign  core_ibuf_io_inst_0_bits_replay = core_ibuf_replay ; 
  assign  core_ibuf_io_inst_0_bits_rvc = core_ibuf__exp_io_rvc ; 
  assign  core_ibuf_io_inst_0_bits_raw = core_ibuf_inst ;
    assign core_ibuf_clock = core_clock;
    assign core_ibuf_reset = core_reset;
    assign core_io_imem_resp_ready = core_ibuf_io_imem_ready;
    assign core_ibuf_io_imem_valid = core_io_imem_resp_valid;
    assign core_ibuf_io_imem_bits_btb_cfiType = core_io_imem_resp_bits_btb_cfiType;
    assign core_ibuf_io_imem_bits_btb_taken = core_io_imem_resp_bits_btb_taken;
    assign core_ibuf_io_imem_bits_btb_mask = core_io_imem_resp_bits_btb_mask;
    assign core_ibuf_io_imem_bits_btb_bridx = core_io_imem_resp_bits_btb_bridx;
    assign core_ibuf_io_imem_bits_btb_target = core_io_imem_resp_bits_btb_target;
    assign core_ibuf_io_imem_bits_btb_entry = core_io_imem_resp_bits_btb_entry;
    assign core_ibuf_io_imem_bits_btb_bht_history = core_io_imem_resp_bits_btb_bht_history;
    assign core_ibuf_io_imem_bits_btb_bht_value = core_io_imem_resp_bits_btb_bht_value;
    assign core_ibuf_io_imem_bits_pc = core_io_imem_resp_bits_pc;
    assign core_ibuf_io_imem_bits_data = core_io_imem_resp_bits_data;
    assign core_ibuf_io_imem_bits_mask = core_io_imem_resp_bits_mask;
    assign core_ibuf_io_imem_bits_xcpt_pf_inst = core_io_imem_resp_bits_xcpt_pf_inst;
    assign core_ibuf_io_imem_bits_xcpt_gf_inst = core_io_imem_resp_bits_xcpt_gf_inst;
    assign core_ibuf_io_imem_bits_xcpt_ae_inst = core_io_imem_resp_bits_xcpt_ae_inst;
    assign core_ibuf_io_imem_bits_replay = core_io_imem_resp_bits_replay;
    assign core_ibuf_io_kill = core_take_pc_mem_wb;
    assign core__ibuf_io_pc = core_ibuf_io_pc;
    assign core__ibuf_io_btb_resp_cfiType = core_ibuf_io_btb_resp_cfiType;
    assign core__ibuf_io_btb_resp_taken = core_ibuf_io_btb_resp_taken;
    assign core__ibuf_io_btb_resp_mask = core_ibuf_io_btb_resp_mask;
    assign core__ibuf_io_btb_resp_bridx = core_ibuf_io_btb_resp_bridx;
    assign core__ibuf_io_btb_resp_target = core_ibuf_io_btb_resp_target;
    assign core__ibuf_io_btb_resp_entry = core_ibuf_io_btb_resp_entry;
    assign core__ibuf_io_btb_resp_bht_history = core_ibuf_io_btb_resp_bht_history;
    assign core__ibuf_io_btb_resp_bht_value = core_ibuf_io_btb_resp_bht_value;
    assign core_ibuf_io_inst_0_ready = ~core_ctrl_stalld;
    assign core__ibuf_io_inst_0_valid = core_ibuf_io_inst_0_valid;
    assign core__ibuf_io_inst_0_bits_xcpt0_pf_inst = core_ibuf_io_inst_0_bits_xcpt0_pf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt0_gf_inst = core_ibuf_io_inst_0_bits_xcpt0_gf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt0_ae_inst = core_ibuf_io_inst_0_bits_xcpt0_ae_inst;
    assign core__ibuf_io_inst_0_bits_xcpt1_pf_inst = core_ibuf_io_inst_0_bits_xcpt1_pf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt1_gf_inst = core_ibuf_io_inst_0_bits_xcpt1_gf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt1_ae_inst = core_ibuf_io_inst_0_bits_xcpt1_ae_inst;
    assign core__ibuf_io_inst_0_bits_replay = core_ibuf_io_inst_0_bits_replay;
    assign core__ibuf_io_inst_0_bits_rvc = core_ibuf_io_inst_0_bits_rvc;
    assign core__ibuf_io_inst_0_bits_inst_bits = core_ibuf_io_inst_0_bits_inst_bits;
    assign core_id_waddr = core_ibuf_io_inst_0_bits_inst_rd;
    assign core__ibuf_io_inst_0_bits_inst_rs1 = core_ibuf_io_inst_0_bits_inst_rs1;
    assign core_id_raddr2 = core_ibuf_io_inst_0_bits_inst_rs2;
    assign core_id_raddr3 = core_ibuf_io_inst_0_bits_inst_rs3;
    assign core__ibuf_io_inst_0_bits_raw = core_ibuf_io_inst_0_bits_raw;
     
  assign  core_id_ctrl_decoder_decoded_plaInput = core__ibuf_io_inst_0_bits_inst_bits ; 
  assign  core_id_raddr1 = core__ibuf_io_inst_0_bits_inst_rs1 ;  
    wire[4:0] core_rf_ext_R0_addr;
    wire core_rf_ext_R0_en;
    wire core_rf_ext_R0_clk;
    wire[31:0] core_rf_ext_R0_data;
    wire[4:0] core_rf_ext_R1_addr;
    wire core_rf_ext_R1_en;
    wire core_rf_ext_R1_clk;
    wire[31:0] core_rf_ext_R1_data;
    wire[4:0] core_rf_ext_W0_addr;
    wire core_rf_ext_W0_en;
    wire core_rf_ext_W0_clk;
    wire[31:0] core_rf_ext_W0_data;

    reg[31:0] core_rf_ext_Memory [0:30]; 
  always @( posedge  core_rf_ext_W0_clk )
         begin 
             if ( core_rf_ext_W0_en &1'h1) 
                 core_rf_ext_Memory  [ core_rf_ext_W0_addr ]<= core_rf_ext_W0_data ;
         end
  assign  core_rf_ext_R0_data = core_rf_ext_R0_en  ?  core_rf_ext_Memory [ core_rf_ext_R0_addr ]:32'bx; 
  assign  core_rf_ext_R1_data = core_rf_ext_R1_en  ?  core_rf_ext_Memory [ core_rf_ext_R1_addr ]:32'bx;
    assign core_rf_ext_R0_addr = ~core_id_raddr2;
    assign core_rf_ext_R0_en = 1'h1;
    assign core_rf_ext_R0_clk = core_clock;
    assign core__rf_ext_R0_data = core_rf_ext_R0_data;
    assign core_rf_ext_R1_addr = ~core_id_raddr1;
    assign core_rf_ext_R1_en = 1'h1;
    assign core_rf_ext_R1_clk = core_clock;
    assign core__rf_ext_R1_data = core_rf_ext_R1_data;
    assign core_rf_ext_W0_addr = ~core_rf_waddr;
    assign core_rf_ext_W0_en = core_rf_wen&(|core_rf_waddr);
    assign core_rf_ext_W0_clk = core_clock;
    assign core_rf_ext_W0_data = core_rf_wdata;
      
    wire core_csr_clock;
    wire core_csr_reset;
    wire core_csr_io_ungated_clock;
    wire core_csr_io_interrupts_debug;
    wire core_csr_io_interrupts_mtip;
    wire core_csr_io_interrupts_msip;
    wire core_csr_io_interrupts_meip;
    wire core_csr_io_hartid;
    wire[11:0] core_csr_io_rw_addr;
    wire[2:0] core_csr_io_rw_cmd;
    wire[31:0] core_csr_io_rw_rdata;
    wire[31:0] core_csr_io_rw_wdata;
    wire[31:0] core_csr_io_decode_0_inst;
    wire core_csr_io_decode_0_read_illegal;
    wire core_csr_io_decode_0_write_illegal;
    wire core_csr_io_decode_0_write_flush;
    wire core_csr_io_decode_0_system_illegal;
    wire core_csr_io_decode_0_virtual_access_illegal;
    wire core_csr_io_decode_0_virtual_system_illegal;
    wire core_csr_io_csr_stall;
    wire core_csr_io_eret;
    wire core_csr_io_singleStep;
    wire core_csr_io_status_debug;
    wire core_csr_io_status_wfi;
    wire[31:0] core_csr_io_status_isa;
    wire core_csr_io_status_dv;
    wire core_csr_io_status_v;
    wire[31:0] core_csr_io_evec;
    wire core_csr_io_exception;
    wire core_csr_io_retire;
    wire[31:0] core_csr_io_cause;
    wire[31:0] core_csr_io_pc;
    wire[31:0] core_csr_io_tval;
    wire[31:0] core_csr_io_htval;
    wire core_csr_io_gva;
    wire[31:0] core_csr_io_time;
    wire core_csr_io_interrupt;
    wire[31:0] core_csr_io_interrupt_cause;
    wire core_csr_io_bp_0_control_action;
    wire[1:0] core_csr_io_bp_0_control_tmatch;
    wire core_csr_io_bp_0_control_x;
    wire core_csr_io_bp_0_control_w;
    wire core_csr_io_bp_0_control_r;
    wire[31:0] core_csr_io_bp_0_address;
    wire core_csr_io_pmp_0_cfg_l;
    wire[1:0] core_csr_io_pmp_0_cfg_a;
    wire core_csr_io_pmp_0_cfg_x;
    wire core_csr_io_pmp_0_cfg_w;
    wire core_csr_io_pmp_0_cfg_r;
    wire[29:0] core_csr_io_pmp_0_addr;
    wire[31:0] core_csr_io_pmp_0_mask;
    wire core_csr_io_pmp_1_cfg_l;
    wire[1:0] core_csr_io_pmp_1_cfg_a;
    wire core_csr_io_pmp_1_cfg_x;
    wire core_csr_io_pmp_1_cfg_w;
    wire core_csr_io_pmp_1_cfg_r;
    wire[29:0] core_csr_io_pmp_1_addr;
    wire[31:0] core_csr_io_pmp_1_mask;
    wire core_csr_io_pmp_2_cfg_l;
    wire[1:0] core_csr_io_pmp_2_cfg_a;
    wire core_csr_io_pmp_2_cfg_x;
    wire core_csr_io_pmp_2_cfg_w;
    wire core_csr_io_pmp_2_cfg_r;
    wire[29:0] core_csr_io_pmp_2_addr;
    wire[31:0] core_csr_io_pmp_2_mask;
    wire core_csr_io_pmp_3_cfg_l;
    wire[1:0] core_csr_io_pmp_3_cfg_a;
    wire core_csr_io_pmp_3_cfg_x;
    wire core_csr_io_pmp_3_cfg_w;
    wire core_csr_io_pmp_3_cfg_r;
    wire[29:0] core_csr_io_pmp_3_addr;
    wire[31:0] core_csr_io_pmp_3_mask;
    wire core_csr_io_pmp_4_cfg_l;
    wire[1:0] core_csr_io_pmp_4_cfg_a;
    wire core_csr_io_pmp_4_cfg_x;
    wire core_csr_io_pmp_4_cfg_w;
    wire core_csr_io_pmp_4_cfg_r;
    wire[29:0] core_csr_io_pmp_4_addr;
    wire[31:0] core_csr_io_pmp_4_mask;
    wire core_csr_io_pmp_5_cfg_l;
    wire[1:0] core_csr_io_pmp_5_cfg_a;
    wire core_csr_io_pmp_5_cfg_x;
    wire core_csr_io_pmp_5_cfg_w;
    wire core_csr_io_pmp_5_cfg_r;
    wire[29:0] core_csr_io_pmp_5_addr;
    wire[31:0] core_csr_io_pmp_5_mask;
    wire core_csr_io_pmp_6_cfg_l;
    wire[1:0] core_csr_io_pmp_6_cfg_a;
    wire core_csr_io_pmp_6_cfg_x;
    wire core_csr_io_pmp_6_cfg_w;
    wire core_csr_io_pmp_6_cfg_r;
    wire[29:0] core_csr_io_pmp_6_addr;
    wire[31:0] core_csr_io_pmp_6_mask;
    wire core_csr_io_pmp_7_cfg_l;
    wire[1:0] core_csr_io_pmp_7_cfg_a;
    wire core_csr_io_pmp_7_cfg_x;
    wire core_csr_io_pmp_7_cfg_w;
    wire core_csr_io_pmp_7_cfg_r;
    wire[29:0] core_csr_io_pmp_7_addr;
    wire[31:0] core_csr_io_pmp_7_mask;
    wire core_csr_io_inhibit_cycle;
    wire[31:0] core_csr_io_inst_0;
    wire core_csr_io_trace_0_valid;
    wire[31:0] core_csr_io_trace_0_iaddr;
    wire[31:0] core_csr_io_trace_0_insn;
    wire[2:0] core_csr_io_trace_0_priv;
    wire core_csr_io_trace_0_exception;
    wire core_csr_io_trace_0_interrupt;
    wire[31:0] core_csr_io_trace_0_cause;
    wire[31:0] core_csr_io_trace_0_tval;
    wire[31:0] core_csr_io_customCSRs_0_value;

    wire[31:0] core_csr__io_rw_rdata_output ; 
    reg core_csr_io_status_cease_r ; 
    wire core_csr__io_csr_stall_output ; 
    wire core_csr__io_singleStep_output ; 
    wire core_csr_mip_meip = core_csr_io_interrupts_meip ; 
    wire core_csr_mip_mtip = core_csr_io_interrupts_mtip ; 
    wire core_csr_mip_msip = core_csr_io_interrupts_msip ; 
    wire[31:0] core_csr_decoded_plaInput_1 = core_csr_io_decode_0_inst ; 
    wire core_csr_reset_mstatus_debug =1'h0; 
    wire core_csr_reset_mstatus_cease =1'h0; 
    wire core_csr_reset_mstatus_wfi =1'h0; 
    wire core_csr_reset_mstatus_dv =1'h0; 
    wire core_csr_reset_mstatus_v =1'h0; 
    wire core_csr_reset_mstatus_sd =1'h0; 
    wire core_csr_reset_mstatus_mpv =1'h0; 
    wire core_csr_reset_mstatus_gva =1'h0; 
    wire core_csr_reset_mstatus_mbe =1'h0; 
    wire core_csr_reset_mstatus_sbe =1'h0; 
    wire core_csr_reset_mstatus_sd_rv32 =1'h0; 
    wire core_csr_reset_mstatus_tsr =1'h0; 
    wire core_csr_reset_mstatus_tw =1'h0; 
    wire core_csr_reset_mstatus_tvm =1'h0; 
    wire core_csr_reset_mstatus_mxr =1'h0; 
    wire core_csr_reset_mstatus_sum =1'h0; 
    wire core_csr_reset_mstatus_mprv =1'h0; 
    wire core_csr_reset_mstatus_spp =1'h0; 
    wire core_csr_reset_mstatus_mpie =1'h0; 
    wire core_csr_reset_mstatus_ube =1'h0; 
    wire core_csr_reset_mstatus_spie =1'h0; 
    wire core_csr_reset_mstatus_upie =1'h0; 
    wire core_csr_reset_mstatus_mie =1'h0; 
    wire core_csr_reset_mstatus_hie =1'h0; 
    wire core_csr_reset_mstatus_sie =1'h0; 
    wire core_csr_reset_mstatus_uie =1'h0; 
    wire core_csr_reset_dcsr_ebreakm =1'h0; 
    wire core_csr_reset_dcsr_ebreakh =1'h0; 
    wire core_csr_reset_dcsr_ebreaks =1'h0; 
    wire core_csr_reset_dcsr_ebreaku =1'h0; 
    wire core_csr_reset_dcsr_zero2 =1'h0; 
    wire core_csr_reset_dcsr_stopcycle =1'h0; 
    wire core_csr_reset_dcsr_stoptime =1'h0; 
    wire core_csr_reset_dcsr_v =1'h0; 
    wire core_csr_reset_dcsr_step =1'h0; 
    wire core_csr_sup_zero1 =1'h0; 
    wire core_csr_sup_debug =1'h0; 
    wire core_csr_sup_rocc =1'h0; 
    wire core_csr_sup_sgeip =1'h0; 
    wire core_csr_sup_vseip =1'h0; 
    wire core_csr_sup_seip =1'h0; 
    wire core_csr_sup_ueip =1'h0; 
    wire core_csr_sup_vstip =1'h0; 
    wire core_csr_sup_stip =1'h0; 
    wire core_csr_sup_utip =1'h0; 
    wire core_csr_sup_vssip =1'h0; 
    wire core_csr_sup_ssip =1'h0; 
    wire core_csr_sup_usip =1'h0; 
    wire core_csr_del_zero1 =1'h0; 
    wire core_csr_del_debug =1'h0; 
    wire core_csr_del_rocc =1'h0; 
    wire core_csr_del_sgeip =1'h0; 
    wire core_csr_del_meip =1'h0; 
    wire core_csr_del_vseip =1'h0; 
    wire core_csr_del_seip =1'h0; 
    wire core_csr_del_ueip =1'h0; 
    wire core_csr_del_mtip =1'h0; 
    wire core_csr_del_vstip =1'h0; 
    wire core_csr_del_stip =1'h0; 
    wire core_csr_del_utip =1'h0; 
    wire core_csr_del_msip =1'h0; 
    wire core_csr_del_vssip =1'h0; 
    wire core_csr_del_ssip =1'h0; 
    wire core_csr_del_usip =1'h0; 
    wire core_csr_always_zero1 =1'h0; 
    wire core_csr_always_debug =1'h0; 
    wire core_csr_always_rocc =1'h0; 
    wire core_csr_always_sgeip =1'h0; 
    wire core_csr_always_meip =1'h0; 
    wire core_csr_always_vseip =1'h0; 
    wire core_csr_always_seip =1'h0; 
    wire core_csr_always_ueip =1'h0; 
    wire core_csr_always_mtip =1'h0; 
    wire core_csr_always_vstip =1'h0; 
    wire core_csr_always_stip =1'h0; 
    wire core_csr_always_utip =1'h0; 
    wire core_csr_always_msip =1'h0; 
    wire core_csr_always_vssip =1'h0; 
    wire core_csr_always_ssip =1'h0; 
    wire core_csr_always_usip =1'h0; 
    wire core_csr_deleg_zero1 =1'h0; 
    wire core_csr_deleg_debug =1'h0; 
    wire core_csr_deleg_rocc =1'h0; 
    wire core_csr_deleg_sgeip =1'h0; 
    wire core_csr_deleg_meip =1'h0; 
    wire core_csr_deleg_vseip =1'h0; 
    wire core_csr_deleg_seip =1'h0; 
    wire core_csr_deleg_ueip =1'h0; 
    wire core_csr_deleg_mtip =1'h0; 
    wire core_csr_deleg_vstip =1'h0; 
    wire core_csr_deleg_stip =1'h0; 
    wire core_csr_deleg_utip =1'h0; 
    wire core_csr_deleg_msip =1'h0; 
    wire core_csr_deleg_vssip =1'h0; 
    wire core_csr_deleg_ssip =1'h0; 
    wire core_csr_deleg_usip =1'h0; 
    wire core_csr_reset_mnstatus_mpv =1'h0; 
    wire core_csr_reset_mnstatus_mie =1'h0; 
    wire core_csr_mip_zero1 =1'h0; 
    wire core_csr_mip_debug =1'h0; 
    wire core_csr_mip_rocc =1'h0; 
    wire core_csr_mip_sgeip =1'h0; 
    wire core_csr_mip_vseip =1'h0; 
    wire core_csr_mip_seip =1'h0; 
    wire core_csr_mip_ueip =1'h0; 
    wire core_csr_mip_vstip =1'h0; 
    wire core_csr_mip_stip =1'h0; 
    wire core_csr_mip_utip =1'h0; 
    wire core_csr_mip_vssip =1'h0; 
    wire core_csr_mip_ssip =1'h0; 
    wire core_csr_mip_usip =1'h0; 
    wire core_csr_lo_hi_5 =1'h0; 
    wire core_csr_hi_hi_5 =1'h0; 
    wire core_csr_read_mnstatus_mpv =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_zero1 =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_debug =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_rocc =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_meip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_vseip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_seip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_ueip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_mtip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_vstip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_stip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_utip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_msip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_vssip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_ssip =1'h0; 
    wire core_csr_sie_mask_sgeip_mask_usip =1'h0; 
    wire core_csr_read_pmp_15_cfg_l =1'h0; 
    wire core_csr_read_pmp_15_cfg_x =1'h0; 
    wire core_csr_read_pmp_15_cfg_w =1'h0; 
    wire core_csr_read_pmp_15_cfg_r =1'h0; 
    wire core_csr_io_decode_0_fp_csr_plaOutput =1'h0; 
    wire core_csr_io_decode_0_read_illegal_plaOutput_1 =1'h0; 
    wire core_csr_delegate =1'h0; 
    wire core_csr_delegateVS =1'h0; 
    wire core_csr_trapToNmiInt =1'h0; 
    wire core_csr_trapToNmiXcpt =1'h0; 
    wire core_csr_trapToNmi =1'h0; 
    wire core_csr_en =1'h0; 
    wire core_csr_delegable =1'h0; 
    wire core_csr_en_1 =1'h0; 
    wire core_csr_delegable_1 =1'h0; 
    wire core_csr_en_2 =1'h0; 
    wire core_csr_delegable_2 =1'h0; 
    wire core_csr_delegable_3 =1'h0; 
    wire core_csr_en_4 =1'h0; 
    wire core_csr_delegable_4 =1'h0; 
    wire core_csr_en_5 =1'h0; 
    wire core_csr_delegable_5 =1'h0; 
    wire core_csr_en_6 =1'h0; 
    wire core_csr_delegable_6 =1'h0; 
    wire core_csr_delegable_7 =1'h0; 
    wire core_csr_en_8 =1'h0; 
    wire core_csr_delegable_8 =1'h0; 
    wire core_csr_en_9 =1'h0; 
    wire core_csr_delegable_9 =1'h0; 
    wire core_csr_en_10 =1'h0; 
    wire core_csr_delegable_10 =1'h0; 
    wire core_csr_delegable_11 =1'h0; 
    wire core_csr_en_12 =1'h0; 
    wire core_csr_delegable_12 =1'h0; 
    wire core_csr_en_13 =1'h0; 
    wire core_csr_delegable_13 =1'h0; 
    wire core_csr_en_14 =1'h0; 
    wire core_csr_delegable_14 =1'h0; 
    wire core_csr_en_15 =1'h0; 
    wire core_csr_delegable_15 =1'h0; 
    wire core_csr_delegable_17 =1'h0; 
    wire core_csr_delegable_21 =1'h0; 
    wire core_csr_delegable_23 =1'h0; 
    wire core_csr_delegable_24 =1'h0; 
    wire core_csr_set_vs_dirty =1'h0; 
    wire core_csr_set_fs_dirty =1'h0; 
    wire core_csr_new_mstatus_debug =1'h0; 
    wire core_csr_new_mstatus_cease =1'h0; 
    wire core_csr_new_mstatus_wfi =1'h0; 
    wire core_csr_new_mstatus_dv =1'h0; 
    wire core_csr_new_mstatus_v =1'h0; 
    wire core_csr_new_mstatus_sd =1'h0; 
    wire core_csr_new_mstatus_mpv =1'h0; 
    wire core_csr_new_mstatus_gva =1'h0; 
    wire core_csr_new_mstatus_mbe =1'h0; 
    wire core_csr_new_mstatus_sbe =1'h0; 
    wire[31:0] core_csr_reset_mstatus_isa =32'h0; 
    wire[31:0] core_csr_read_mideleg =32'h0; 
    wire[31:0] core_csr_read_medeleg =32'h0; 
    wire[31:0] core_csr_read_mcounteren =32'h0; 
    wire[31:0] core_csr_read_scounteren =32'h0; 
    wire[31:0] core_csr_read_hideleg =32'h0; 
    wire[31:0] core_csr_read_hedeleg =32'h0; 
    wire[31:0] core_csr_read_hcounteren =32'h0; 
    wire[31:0] core_csr_read_hie =32'h0; 
    wire[31:0] core_csr_read_vstvec =32'h0; 
    wire[31:0] core_csr_s_interrupts =32'h0; 
    wire[31:0] core_csr_vs_interrupts =32'h0; 
    wire[31:0] core_csr_read_stvec =32'h0; 
    wire[31:0] core_csr_sie_mask =32'h0; 
    wire[31:0] core_csr_read_pmp_15_mask =32'h0; 
    wire[31:0] core_csr_new_mstatus_isa =32'h0; 
    wire[15:0] core_csr_delegable_interrupts =16'h0; 
    wire[15:0] core_csr_hs_delegable_interrupts =16'h0; 
    wire[15:0] core_csr_mideleg_always_hs =16'h0; 
    wire[15:0] core_csr_read_hvip =16'h0; 
    wire[15:0] core_csr_read_hip =16'h0; 
    wire[15:0] core_csr_lo_21 =16'h0; 
    wire[15:0] core_csr_hi_21 =16'h0; 
    wire[15:0] core_csr_lo_26 =16'h0; 
    wire[15:0] core_csr_hi_26 =16'h0; 
    wire[3:0] core_csr_hi_hi =4'h0; 
    wire[3:0] core_csr_lo_lo_1 =4'h0; 
    wire[3:0] core_csr_lo_hi_1 =4'h0; 
    wire[3:0] core_csr_hi_lo_1 =4'h0; 
    wire[3:0] core_csr_hi_hi_1 =4'h0; 
    wire[3:0] core_csr_lo_lo_2 =4'h0; 
    wire[3:0] core_csr_lo_hi_2 =4'h0; 
    wire[3:0] core_csr_hi_lo_2 =4'h0; 
    wire[3:0] core_csr_hi_hi_2 =4'h0; 
    wire[3:0] core_csr_lo_lo_3 =4'h0; 
    wire[3:0] core_csr_lo_hi_3 =4'h0; 
    wire[3:0] core_csr_hi_lo_3 =4'h0; 
    wire[3:0] core_csr_hi_hi_3 =4'h0; 
    wire[3:0] core_csr_read_mstatus_lo_hi_lo_hi =4'h0; 
    wire[3:0] core_csr_hi_lo_5 =4'h0; 
    wire[3:0] core_csr_sie_mask_lo_lo =4'h0; 
    wire[3:0] core_csr_sie_mask_lo_hi =4'h0; 
    wire[3:0] core_csr_sie_mask_hi_lo =4'h0; 
    wire[3:0] core_csr_decoded_orMatrixOutputs_lo =4'h0; 
    wire[3:0] core_csr_decoded_orMatrixOutputs_lo_1 =4'h0; 
    wire[3:0] core_csr_newBPC_lo_hi_1 =4'h0; 
    wire[3:0] core_csr_newBPC_hi_lo_lo_1 =4'h0; 
    wire[2:0] core_csr_reset_dcsr_cause =3'h0; 
    wire[2:0] core_csr_reset_mnstatus_zero3 =3'h0; 
    wire[2:0] core_csr_reset_mnstatus_zero2 =3'h0; 
    wire[2:0] core_csr_reset_mnstatus_zero1 =3'h0; 
    wire[2:0] core_csr_read_mstatus_lo_hi_hi_hi =3'h0; 
    wire[2:0] core_csr_read_mstatus_hi_lo_lo_hi =3'h0; 
    wire[2:0] core_csr_read_mstatus_hi_lo_hi_lo =3'h0; 
    wire[2:0] core_csr_read_mnstatus_zero3 =3'h0; 
    wire[2:0] core_csr_read_mnstatus_zero2 =3'h0; 
    wire[2:0] core_csr_read_mnstatus_zero1 =3'h0; 
    wire[2:0] core_csr_lo_17 =3'h0; 
    wire[2:0] core_csr_hi_hi_15 =3'h0; 
    wire[2:0] core_csr_lo_18 =3'h0; 
    wire[2:0] core_csr_hi_hi_16 =3'h0; 
    wire[2:0] core_csr_lo_19 =3'h0; 
    wire[2:0] core_csr_hi_hi_17 =3'h0; 
    wire[2:0] core_csr_lo_20 =3'h0; 
    wire[2:0] core_csr_hi_hi_18 =3'h0; 
    wire[2:0] core_csr_lo_22 =3'h0; 
    wire[2:0] core_csr_hi_hi_19 =3'h0; 
    wire[2:0] core_csr_lo_23 =3'h0; 
    wire[2:0] core_csr_hi_hi_20 =3'h0; 
    wire[2:0] core_csr_lo_24 =3'h0; 
    wire[2:0] core_csr_hi_hi_21 =3'h0; 
    wire[2:0] core_csr_lo_25 =3'h0; 
    wire[2:0] core_csr_hi_hi_22 =3'h0; 
    wire[2:0] core_csr_newBPC_lo_lo_1 =3'h0; 
    wire[1:0] core_csr_reset_mstatus_dprv =2'h0; 
    wire[1:0] core_csr_reset_mstatus_sxl =2'h0; 
    wire[1:0] core_csr_reset_mstatus_uxl =2'h0; 
    wire[1:0] core_csr_reset_mstatus_xs =2'h0; 
    wire[1:0] core_csr_reset_mstatus_fs =2'h0; 
    wire[1:0] core_csr_reset_mstatus_vs =2'h0; 
    wire[1:0] core_csr_reset_dcsr_zero4 =2'h0; 
    wire[1:0] core_csr_reset_dcsr_zero1 =2'h0; 
    wire[1:0] core_csr_lo_lo_lo =2'h0; 
    wire[1:0] core_csr_lo_hi_lo =2'h0; 
    wire[1:0] core_csr_hi_lo_lo =2'h0; 
    wire[1:0] core_csr_hi_hi_lo =2'h0; 
    wire[1:0] core_csr_hi_hi_hi =2'h0; 
    wire[1:0] core_csr_lo_lo_lo_1 =2'h0; 
    wire[1:0] core_csr_lo_lo_hi_1 =2'h0; 
    wire[1:0] core_csr_lo_hi_lo_1 =2'h0; 
    wire[1:0] core_csr_lo_hi_hi_1 =2'h0; 
    wire[1:0] core_csr_hi_lo_lo_1 =2'h0; 
    wire[1:0] core_csr_hi_lo_hi_1 =2'h0; 
    wire[1:0] core_csr_hi_hi_lo_1 =2'h0; 
    wire[1:0] core_csr_hi_hi_hi_1 =2'h0; 
    wire[1:0] core_csr_lo_lo_lo_2 =2'h0; 
    wire[1:0] core_csr_lo_lo_hi_2 =2'h0; 
    wire[1:0] core_csr_lo_hi_lo_2 =2'h0; 
    wire[1:0] core_csr_lo_hi_hi_2 =2'h0; 
    wire[1:0] core_csr_hi_lo_lo_2 =2'h0; 
    wire[1:0] core_csr_hi_lo_hi_2 =2'h0; 
    wire[1:0] core_csr_hi_hi_lo_2 =2'h0; 
    wire[1:0] core_csr_hi_hi_hi_2 =2'h0; 
    wire[1:0] core_csr_lo_lo_lo_3 =2'h0; 
    wire[1:0] core_csr_lo_lo_hi_3 =2'h0; 
    wire[1:0] core_csr_lo_hi_lo_3 =2'h0; 
    wire[1:0] core_csr_lo_hi_hi_3 =2'h0; 
    wire[1:0] core_csr_hi_lo_lo_3 =2'h0; 
    wire[1:0] core_csr_hi_lo_hi_3 =2'h0; 
    wire[1:0] core_csr_hi_hi_lo_3 =2'h0; 
    wire[1:0] core_csr_hi_hi_hi_3 =2'h0; 
    wire[1:0] core_csr_read_hvip_lo_lo_lo =2'h0; 
    wire[1:0] core_csr_read_hvip_lo_lo_hi =2'h0; 
    wire[1:0] core_csr_read_hvip_lo_hi_lo =2'h0; 
    wire[1:0] core_csr_read_hvip_lo_hi_hi =2'h0; 
    wire[1:0] core_csr_read_hvip_hi_lo_lo =2'h0; 
    wire[1:0] core_csr_read_hvip_hi_lo_hi =2'h0; 
    wire[1:0] core_csr_read_hvip_hi_hi_lo =2'h0; 
    wire[1:0] core_csr_read_hvip_hi_hi_hi =2'h0; 
    wire[1:0] core_csr_pmp_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_1_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_2_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_3_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_4_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_5_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_6_cfg_res =2'h0; 
    wire[1:0] core_csr_pmp_7_cfg_res =2'h0; 
    wire[1:0] core_csr_read_mstatus_lo_lo_lo_lo =2'h0; 
    wire[1:0] core_csr_read_mstatus_lo_lo_hi_lo =2'h0; 
    wire[1:0] core_csr_read_mstatus_lo_hi_hi_lo =2'h0; 
    wire[1:0] core_csr_read_mstatus_lo_hi_hi_hi_hi =2'h0; 
    wire[1:0] core_csr_lo_hi_lo_4 =2'h0; 
    wire[1:0] core_csr_lo_hi_hi_5 =2'h0; 
    wire[1:0] core_csr_hi_lo_lo_5 =2'h0; 
    wire[1:0] core_csr_hi_lo_hi_5 =2'h0; 
    wire[1:0] core_csr_read_vcsr =2'h0; 
    wire[1:0] core_csr_sie_mask_lo_lo_lo =2'h0; 
    wire[1:0] core_csr_sie_mask_lo_lo_hi =2'h0; 
    wire[1:0] core_csr_sie_mask_lo_hi_lo =2'h0; 
    wire[1:0] core_csr_sie_mask_lo_hi_hi =2'h0; 
    wire[1:0] core_csr_sie_mask_hi_lo_lo =2'h0; 
    wire[1:0] core_csr_sie_mask_hi_lo_hi =2'h0; 
    wire[1:0] core_csr_sie_mask_hi_hi_hi =2'h0; 
    wire[1:0] core_csr_read_pmp_15_cfg_res =2'h0; 
    wire[1:0] core_csr_read_pmp_15_cfg_a =2'h0; 
    wire[1:0] core_csr_lo_hi_15 =2'h0; 
    wire[1:0] core_csr_lo_hi_16 =2'h0; 
    wire[1:0] core_csr_lo_hi_17 =2'h0; 
    wire[1:0] core_csr_lo_hi_18 =2'h0; 
    wire[1:0] core_csr_lo_hi_19 =2'h0; 
    wire[1:0] core_csr_lo_hi_20 =2'h0; 
    wire[1:0] core_csr_lo_hi_21 =2'h0; 
    wire[1:0] core_csr_lo_hi_22 =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_lo =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_hi =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_lo_1 =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_hi_1 =2'h0; 
    wire[1:0] core_csr_causeIsDebugBreak_lo =2'h0; 
    wire[1:0] core_csr_nmiTVec =2'h0; 
    wire[1:0] core_csr_new_mstatus_dprv =2'h0; 
    wire[1:0] core_csr_new_mstatus_prv =2'h0; 
    wire[1:0] core_csr_new_mstatus_sxl =2'h0; 
    wire[1:0] core_csr_new_mstatus_uxl =2'h0; 
    wire[1:0] core_csr_new_mip_lo_lo_lo =2'h0; 
    wire[1:0] core_csr_new_mip_lo_lo_hi =2'h0; 
    wire[1:0] core_csr_new_mip_lo_hi_lo =2'h0; 
    wire[1:0] core_csr_new_mip_lo_hi_hi =2'h0; 
    wire[1:0] core_csr_new_mip_hi_lo_lo =2'h0; 
    wire[1:0] core_csr_new_mip_hi_lo_hi =2'h0; 
    wire[1:0] core_csr_new_mip_hi_hi_lo =2'h0; 
    wire[1:0] core_csr_new_mip_hi_hi_hi =2'h0; 
    wire[1:0] core_csr_newBPC_lo_hi_lo =2'h0; 
    wire[1:0] core_csr_newBPC_lo_lo_hi_1 =2'h0; 
    wire[1:0] core_csr_newBPC_lo_hi_lo_1 =2'h0; 
    wire[1:0] core_csr_newBPC_lo_hi_hi_1 =2'h0; 
    wire[1:0] core_csr_newBPC_hi_lo_hi_1 =2'h0; 
    wire[22:0] core_csr_reset_mstatus_zero2 =23'h0; 
    wire[22:0] core_csr_new_mstatus_zero2 =23'h0; 
    wire core_csr_sup_meip =1'h1; 
    wire core_csr_sup_mtip =1'h1; 
    wire core_csr_sup_msip =1'h1; 
    wire core_csr_read_mnstatus_mie =1'h1; 
    wire core_csr_sie_mask_sgeip_mask_sgeip =1'h1; 
    wire core_csr_allow_wfi =1'h1; 
    wire core_csr_allow_sfence_vma =1'h1; 
    wire core_csr_allow_hfence_vvma =1'h1; 
    wire core_csr_allow_hlsv =1'h1; 
    wire core_csr_allow_sret =1'h1; 
    wire core_csr_allow_counter =1'h1; 
    wire core_csr_csr_addr_legal =1'h1; 
    wire core_csr_delegable_16 =1'h1; 
    wire core_csr_delegable_18 =1'h1; 
    wire core_csr_delegable_19 =1'h1; 
    wire core_csr_delegable_20 =1'h1; 
    wire core_csr_delegable_22 =1'h1; 
    wire[3:0] core_csr_lo_lo =4'h8; 
    wire[3:0] core_csr_lo_hi =4'h8; 
    wire[3:0] core_csr_hi_lo =4'h8; 
    wire[3:0] core_csr_lo_hi_4 =4'h8; 
    wire[3:0] core_csr_newBPC_lo_hi =4'h8; 
    wire[3:0] core_csr_sie_mask_hi_hi =4'h1; 
    wire[6:0] core_csr_newBPC_lo_1 =7'h0; 
    wire[1:0] core_csr_reset_mstatus_prv =2'h3; 
    wire[1:0] core_csr_reset_mstatus_mpp =2'h3; 
    wire[1:0] core_csr_reset_dcsr_prv =2'h3; 
    wire[1:0] core_csr_reset_mnstatus_mpp =2'h3; 
    wire[1:0] core_csr_read_mnstatus_mpp =2'h3; 
    wire[8:0] core_csr_read_mstatus_hi_lo_lo_lo =9'h0; 
    wire[24:0] core_csr_newBPC_hi_1 =25'h0; 
    wire[18:0] core_csr_newBPC_hi_hi_1 =19'h0; 
    wire[4:0] core_csr_read_mstatus_lo_hi_hi =5'h0; 
    wire[4:0] core_csr_hi_17 =5'h0; 
    wire[4:0] core_csr_hi_18 =5'h0; 
    wire[4:0] core_csr_hi_19 =5'h0; 
    wire[4:0] core_csr_hi_20 =5'h0; 
    wire[4:0] core_csr_hi_22 =5'h0; 
    wire[4:0] core_csr_hi_23 =5'h0; 
    wire[4:0] core_csr_hi_24 =5'h0; 
    wire[4:0] core_csr_hi_25 =5'h0; 
    wire[4:0] core_csr_newBPC_hi_hi_hi_1 =5'h0; 
    wire[13:0] core_csr_newBPC_hi_hi_lo_1 =14'h0; 
    wire[5:0] core_csr_newBPC_hi_lo_1 =6'h0; 
    wire[13:0] core_csr_hi_hi_lo_4 =14'h400; 
    wire[13:0] core_csr_newBPC_hi_hi_lo =14'h400; 
    wire[1:0] core_csr_lo_lo_hi =2'h2; 
    wire[1:0] core_csr_lo_hi_hi =2'h2; 
    wire[1:0] core_csr_hi_lo_hi =2'h2; 
    wire[1:0] core_csr_lo_hi_hi_4 =2'h2; 
    wire[1:0] core_csr_newBPC_lo_hi_hi =2'h2; 
    wire[3:0] core_csr_hi_hi_hi_5 =4'h4; 
    wire[23:0] core_csr_read_mstatus_hi_hi_lo_lo =24'h0; 
    wire[23:0] core_csr_hi_5 =24'h0; 
    wire[11:0] core_csr_reset_dcsr_zero3 =12'h0; 
    wire[11:0] core_csr_read_mstatus_hi_lo_lo =12'h0; 
    wire[7:0] core_csr_reset_mstatus_zero1 =8'h0; 
    wire[7:0] core_csr_lo_1 =8'h0; 
    wire[7:0] core_csr_hi_1 =8'h0; 
    wire[7:0] core_csr_lo_2 =8'h0; 
    wire[7:0] core_csr_hi_2 =8'h0; 
    wire[7:0] core_csr_lo_3 =8'h0; 
    wire[7:0] core_csr_hi_3 =8'h0; 
    wire[7:0] core_csr_read_fcsr =8'h0; 
    wire[7:0] core_csr_sie_mask_lo =8'h0; 
    wire[7:0] core_csr_lo =8'h88; 
    wire[7:0] core_csr_hi =8'h8; 
    wire[15:0] core_csr_supported_interrupts =16'h888; 
    wire[1:0] core_csr_reset_dcsr_xdebugver =2'h1; 
    wire[1:0] core_csr_sie_mask_hi_hi_lo =2'h1; 
    wire[7:0] core_csr_sie_mask_hi =8'h10; 
    wire[29:0] core_csr_read_pmp_15_addr =30'h0; 
    reg core_csr_reg_mstatus_v ; 
    reg core_csr_reg_mstatus_mpv ; 
    reg core_csr_reg_mstatus_gva ; reg[1:0] core_csr_reg_mstatus_mpp ; 
    reg core_csr_reg_mstatus_mpie ; 
    reg core_csr_reg_mstatus_mie ; 
    reg core_csr_reg_dcsr_ebreakm ; reg[2:0] core_csr_reg_dcsr_cause ; 
    reg core_csr_reg_dcsr_v ; 
    reg core_csr_reg_dcsr_step ; 
    reg core_csr_reg_debug ; reg[31:0] core_csr_reg_dpc ; reg[31:0] core_csr_reg_dscratch0 ; 
    reg core_csr_reg_singleStepped ; 
    reg core_csr_reg_bp_0_control_dmode ; 
    reg core_csr_reg_bp_0_control_action ; reg[1:0] core_csr_reg_bp_0_control_tmatch ; 
    reg core_csr_reg_bp_0_control_x ; 
    reg core_csr_reg_bp_0_control_w ; 
    reg core_csr_reg_bp_0_control_r ; reg[31:0] core_csr_reg_bp_0_address ; 
    reg core_csr_reg_pmp_0_cfg_l ; 
    wire core_csr_pmp_cfg_l = core_csr_reg_pmp_0_cfg_l ; reg[1:0] core_csr_reg_pmp_0_cfg_a ; 
    wire[1:0] core_csr_pmp_cfg_a = core_csr_reg_pmp_0_cfg_a ; 
    reg core_csr_reg_pmp_0_cfg_x ; 
    wire core_csr_pmp_cfg_x = core_csr_reg_pmp_0_cfg_x ; 
    reg core_csr_reg_pmp_0_cfg_w ; 
    wire core_csr_pmp_cfg_w = core_csr_reg_pmp_0_cfg_w ; 
    reg core_csr_reg_pmp_0_cfg_r ; 
    wire core_csr_pmp_cfg_r = core_csr_reg_pmp_0_cfg_r ; reg[29:0] core_csr_reg_pmp_0_addr ; 
    wire[29:0] core_csr_pmp_addr = core_csr_reg_pmp_0_addr ; 
    reg core_csr_reg_pmp_1_cfg_l ; 
    wire core_csr_pmp_1_cfg_l = core_csr_reg_pmp_1_cfg_l ; reg[1:0] core_csr_reg_pmp_1_cfg_a ; 
    wire[1:0] core_csr_pmp_1_cfg_a = core_csr_reg_pmp_1_cfg_a ; 
    reg core_csr_reg_pmp_1_cfg_x ; 
    wire core_csr_pmp_1_cfg_x = core_csr_reg_pmp_1_cfg_x ; 
    reg core_csr_reg_pmp_1_cfg_w ; 
    wire core_csr_pmp_1_cfg_w = core_csr_reg_pmp_1_cfg_w ; 
    reg core_csr_reg_pmp_1_cfg_r ; 
    wire core_csr_pmp_1_cfg_r = core_csr_reg_pmp_1_cfg_r ; reg[29:0] core_csr_reg_pmp_1_addr ; 
    wire[29:0] core_csr_pmp_1_addr = core_csr_reg_pmp_1_addr ; 
    reg core_csr_reg_pmp_2_cfg_l ; 
    wire core_csr_pmp_2_cfg_l = core_csr_reg_pmp_2_cfg_l ; reg[1:0] core_csr_reg_pmp_2_cfg_a ; 
    wire[1:0] core_csr_pmp_2_cfg_a = core_csr_reg_pmp_2_cfg_a ; 
    reg core_csr_reg_pmp_2_cfg_x ; 
    wire core_csr_pmp_2_cfg_x = core_csr_reg_pmp_2_cfg_x ; 
    reg core_csr_reg_pmp_2_cfg_w ; 
    wire core_csr_pmp_2_cfg_w = core_csr_reg_pmp_2_cfg_w ; 
    reg core_csr_reg_pmp_2_cfg_r ; 
    wire core_csr_pmp_2_cfg_r = core_csr_reg_pmp_2_cfg_r ; reg[29:0] core_csr_reg_pmp_2_addr ; 
    wire[29:0] core_csr_pmp_2_addr = core_csr_reg_pmp_2_addr ; 
    reg core_csr_reg_pmp_3_cfg_l ; 
    wire core_csr_pmp_3_cfg_l = core_csr_reg_pmp_3_cfg_l ; reg[1:0] core_csr_reg_pmp_3_cfg_a ; 
    wire[1:0] core_csr_pmp_3_cfg_a = core_csr_reg_pmp_3_cfg_a ; 
    reg core_csr_reg_pmp_3_cfg_x ; 
    wire core_csr_pmp_3_cfg_x = core_csr_reg_pmp_3_cfg_x ; 
    reg core_csr_reg_pmp_3_cfg_w ; 
    wire core_csr_pmp_3_cfg_w = core_csr_reg_pmp_3_cfg_w ; 
    reg core_csr_reg_pmp_3_cfg_r ; 
    wire core_csr_pmp_3_cfg_r = core_csr_reg_pmp_3_cfg_r ; reg[29:0] core_csr_reg_pmp_3_addr ; 
    wire[29:0] core_csr_pmp_3_addr = core_csr_reg_pmp_3_addr ; 
    reg core_csr_reg_pmp_4_cfg_l ; 
    wire core_csr_pmp_4_cfg_l = core_csr_reg_pmp_4_cfg_l ; reg[1:0] core_csr_reg_pmp_4_cfg_a ; 
    wire[1:0] core_csr_pmp_4_cfg_a = core_csr_reg_pmp_4_cfg_a ; 
    reg core_csr_reg_pmp_4_cfg_x ; 
    wire core_csr_pmp_4_cfg_x = core_csr_reg_pmp_4_cfg_x ; 
    reg core_csr_reg_pmp_4_cfg_w ; 
    wire core_csr_pmp_4_cfg_w = core_csr_reg_pmp_4_cfg_w ; 
    reg core_csr_reg_pmp_4_cfg_r ; 
    wire core_csr_pmp_4_cfg_r = core_csr_reg_pmp_4_cfg_r ; reg[29:0] core_csr_reg_pmp_4_addr ; 
    wire[29:0] core_csr_pmp_4_addr = core_csr_reg_pmp_4_addr ; 
    reg core_csr_reg_pmp_5_cfg_l ; 
    wire core_csr_pmp_5_cfg_l = core_csr_reg_pmp_5_cfg_l ; reg[1:0] core_csr_reg_pmp_5_cfg_a ; 
    wire[1:0] core_csr_pmp_5_cfg_a = core_csr_reg_pmp_5_cfg_a ; 
    reg core_csr_reg_pmp_5_cfg_x ; 
    wire core_csr_pmp_5_cfg_x = core_csr_reg_pmp_5_cfg_x ; 
    reg core_csr_reg_pmp_5_cfg_w ; 
    wire core_csr_pmp_5_cfg_w = core_csr_reg_pmp_5_cfg_w ; 
    reg core_csr_reg_pmp_5_cfg_r ; 
    wire core_csr_pmp_5_cfg_r = core_csr_reg_pmp_5_cfg_r ; reg[29:0] core_csr_reg_pmp_5_addr ; 
    wire[29:0] core_csr_pmp_5_addr = core_csr_reg_pmp_5_addr ; 
    reg core_csr_reg_pmp_6_cfg_l ; 
    wire core_csr_pmp_6_cfg_l = core_csr_reg_pmp_6_cfg_l ; reg[1:0] core_csr_reg_pmp_6_cfg_a ; 
    wire[1:0] core_csr_pmp_6_cfg_a = core_csr_reg_pmp_6_cfg_a ; 
    reg core_csr_reg_pmp_6_cfg_x ; 
    wire core_csr_pmp_6_cfg_x = core_csr_reg_pmp_6_cfg_x ; 
    reg core_csr_reg_pmp_6_cfg_w ; 
    wire core_csr_pmp_6_cfg_w = core_csr_reg_pmp_6_cfg_w ; 
    reg core_csr_reg_pmp_6_cfg_r ; 
    wire core_csr_pmp_6_cfg_r = core_csr_reg_pmp_6_cfg_r ; reg[29:0] core_csr_reg_pmp_6_addr ; 
    wire[29:0] core_csr_pmp_6_addr = core_csr_reg_pmp_6_addr ; 
    reg core_csr_reg_pmp_7_cfg_l ; 
    wire core_csr_pmp_7_cfg_l = core_csr_reg_pmp_7_cfg_l ; reg[1:0] core_csr_reg_pmp_7_cfg_a ; 
    wire[1:0] core_csr_pmp_7_cfg_a = core_csr_reg_pmp_7_cfg_a ; 
    reg core_csr_reg_pmp_7_cfg_x ; 
    wire core_csr_pmp_7_cfg_x = core_csr_reg_pmp_7_cfg_x ; 
    reg core_csr_reg_pmp_7_cfg_w ; 
    wire core_csr_pmp_7_cfg_w = core_csr_reg_pmp_7_cfg_w ; 
    reg core_csr_reg_pmp_7_cfg_r ; 
    wire core_csr_pmp_7_cfg_r = core_csr_reg_pmp_7_cfg_r ; reg[29:0] core_csr_reg_pmp_7_addr ; 
    wire[29:0] core_csr_pmp_7_addr = core_csr_reg_pmp_7_addr ; reg[31:0] core_csr_reg_mie ; reg[31:0] core_csr_reg_mepc ; reg[31:0] core_csr_reg_mcause ; reg[31:0] core_csr_reg_mtval ; reg[31:0] core_csr_reg_mtval2 ; reg[31:0] core_csr_reg_mscratch ; reg[31:0] core_csr_reg_mtvec ; 
    wire[3:0] core_csr_read_hvip_lo_lo ={ core_csr_read_hvip_lo_lo_hi , core_csr_read_hvip_lo_lo_lo }; 
    wire[3:0] core_csr_read_hvip_lo_hi ={ core_csr_read_hvip_lo_hi_hi , core_csr_read_hvip_lo_hi_lo }; 
    wire[7:0] core_csr_read_hvip_lo ={ core_csr_read_hvip_lo_hi , core_csr_read_hvip_lo_lo }; 
    wire[3:0] core_csr_read_hvip_hi_lo ={ core_csr_read_hvip_hi_lo_hi , core_csr_read_hvip_hi_lo_lo }; 
    wire[3:0] core_csr_read_hvip_hi_hi ={ core_csr_read_hvip_hi_hi_hi , core_csr_read_hvip_hi_hi_lo }; 
    wire[7:0] core_csr_read_hvip_hi ={ core_csr_read_hvip_hi_hi , core_csr_read_hvip_hi_lo }; 
    reg core_csr_reg_wfi ; reg[2:0] core_csr_reg_mcountinhibit ; 
    wire core_csr_x11 = core_csr_reg_mcountinhibit [0]; 
    wire core_csr_x3 = core_csr_reg_mcountinhibit [2]; reg[5:0] core_csr_small_0 ; 
    wire[6:0] core_csr_nextSmall ={1'h0, core_csr_small_0 }+{6'h0, core_csr_io_retire }; reg[57:0] core_csr_large_0 ; 
    wire[63:0] core_csr_value ={ core_csr_large_0 , core_csr_small_0 }; 
    wire core_csr_x10 =~ core_csr__io_csr_stall_output ; reg[5:0] core_csr_small_1 ; 
    wire[6:0] core_csr_nextSmall_1 ={1'h0, core_csr_small_1 }+{6'h0, core_csr_x10 }; reg[57:0] core_csr_large_1 ; 
    wire[63:0] core_csr_value_1 ={ core_csr_large_1 , core_csr_small_1 }; 
    wire[1:0] core_csr_read_mip_lo_lo_lo ={ core_csr_mip_ssip , core_csr_mip_usip }; 
    wire[1:0] core_csr_read_mip_lo_lo_hi ={ core_csr_mip_msip , core_csr_mip_vssip }; 
    wire[3:0] core_csr_read_mip_lo_lo ={ core_csr_read_mip_lo_lo_hi , core_csr_read_mip_lo_lo_lo }; 
    wire[1:0] core_csr_read_mip_lo_hi_lo ={ core_csr_mip_stip , core_csr_mip_utip }; 
    wire[1:0] core_csr_read_mip_lo_hi_hi ={ core_csr_mip_mtip , core_csr_mip_vstip }; 
    wire[3:0] core_csr_read_mip_lo_hi ={ core_csr_read_mip_lo_hi_hi , core_csr_read_mip_lo_hi_lo }; 
    wire[7:0] core_csr_read_mip_lo ={ core_csr_read_mip_lo_hi , core_csr_read_mip_lo_lo }; 
    wire[1:0] core_csr_read_mip_hi_lo_lo ={ core_csr_mip_seip , core_csr_mip_ueip }; 
    wire[1:0] core_csr_read_mip_hi_lo_hi ={ core_csr_mip_meip , core_csr_mip_vseip }; 
    wire[3:0] core_csr_read_mip_hi_lo ={ core_csr_read_mip_hi_lo_hi , core_csr_read_mip_hi_lo_lo }; 
    wire[1:0] core_csr_read_mip_hi_hi_lo ={1'h0, core_csr_mip_sgeip }; 
    wire[1:0] core_csr_read_mip_hi_hi_hi ={ core_csr_mip_zero1 , core_csr_mip_debug }; 
    wire[3:0] core_csr_read_mip_hi_hi ={ core_csr_read_mip_hi_hi_hi , core_csr_read_mip_hi_hi_lo }; 
    wire[7:0] core_csr_read_mip_hi ={ core_csr_read_mip_hi_hi , core_csr_read_mip_hi_lo }; 
    wire[15:0] core_csr_read_mip ={ core_csr_read_mip_hi , core_csr_read_mip_lo }&16'h888; 
    wire[31:0] core_csr_pending_interrupts ={16'h0, core_csr_reg_mie [15:0]& core_csr_read_mip }; 
    wire[14:0] core_csr_d_interrupts ={ core_csr_io_interrupts_debug ,14'h0}; 
    wire[31:0] core_csr_m_interrupts = core_csr_reg_mstatus_mie  ?  core_csr_pending_interrupts :32'h0; 
    wire core_csr_anyInterrupt =(| core_csr_d_interrupts )| core_csr_m_interrupts [15]| core_csr_m_interrupts [14]| core_csr_m_interrupts [13]| core_csr_m_interrupts [12]| core_csr_m_interrupts [11]| core_csr_m_interrupts [3]| core_csr_m_interrupts [7]| core_csr_m_interrupts [9]| core_csr_m_interrupts [1]| core_csr_m_interrupts [5]| core_csr_m_interrupts [10]| core_csr_m_interrupts [2]| core_csr_m_interrupts [6]| core_csr_m_interrupts [8]| core_csr_m_interrupts [0]| core_csr_m_interrupts [4]; 
    wire[3:0] core_csr_whichInterrupt = core_csr_d_interrupts [14] ? 4'hE: core_csr_d_interrupts [13] ? 4'hD: core_csr_d_interrupts [12] ? 4'hC: core_csr_d_interrupts [11] ? 4'hB: core_csr_d_interrupts [3] ? 4'h3: core_csr_d_interrupts [7] ? 4'h7: core_csr_d_interrupts [9] ? 4'h9: core_csr_d_interrupts [1] ? 4'h1: core_csr_d_interrupts [5] ? 4'h5: core_csr_d_interrupts [10] ? 4'hA: core_csr_d_interrupts [2] ? 4'h2: core_csr_d_interrupts [6] ? 4'h6: core_csr_d_interrupts [8] ? 4'h8: core_csr_d_interrupts [0] ? 4'h0: core_csr_d_interrupts [4] ? 4'h4: core_csr_m_interrupts [15] ? 4'hF: core_csr_m_interrupts [14] ? 4'hE: core_csr_m_interrupts [13] ? 4'hD: core_csr_m_interrupts [12] ? 4'hC: core_csr_m_interrupts [11] ? 4'hB: core_csr_m_interrupts [3] ? 4'h3: core_csr_m_interrupts [7] ? 4'h7: core_csr_m_interrupts [9] ? 4'h9: core_csr_m_interrupts [1] ? 4'h1: core_csr_m_interrupts [5] ? 4'h5: core_csr_m_interrupts [10] ? 4'hA: core_csr_m_interrupts [2] ? 4'h2: core_csr_m_interrupts [6] ? 4'h6: core_csr_m_interrupts [8] ? 4'h8:{1'h0,~( core_csr_m_interrupts [0]),2'h0}; 
    wire[31:0] core_csr_interruptCause ={28'h0, core_csr_whichInterrupt }-32'h80000000; 
    wire[30:0] core_csr_pmp_mask_base ={ core_csr_pmp_addr , core_csr_pmp_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_mask ={ core_csr_pmp_mask_base [29:0]&~( core_csr_pmp_mask_base [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_1 ={ core_csr_pmp_1_addr , core_csr_pmp_1_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_1_mask ={ core_csr_pmp_mask_base_1 [29:0]&~( core_csr_pmp_mask_base_1 [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_2 ={ core_csr_pmp_2_addr , core_csr_pmp_2_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_2_mask ={ core_csr_pmp_mask_base_2 [29:0]&~( core_csr_pmp_mask_base_2 [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_3 ={ core_csr_pmp_3_addr , core_csr_pmp_3_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_3_mask ={ core_csr_pmp_mask_base_3 [29:0]&~( core_csr_pmp_mask_base_3 [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_4 ={ core_csr_pmp_4_addr , core_csr_pmp_4_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_4_mask ={ core_csr_pmp_mask_base_4 [29:0]&~( core_csr_pmp_mask_base_4 [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_5 ={ core_csr_pmp_5_addr , core_csr_pmp_5_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_5_mask ={ core_csr_pmp_mask_base_5 [29:0]&~( core_csr_pmp_mask_base_5 [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_6 ={ core_csr_pmp_6_addr , core_csr_pmp_6_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_6_mask ={ core_csr_pmp_mask_base_6 [29:0]&~( core_csr_pmp_mask_base_6 [29:0]+30'h1),2'h3}; 
    wire[30:0] core_csr_pmp_mask_base_7 ={ core_csr_pmp_7_addr , core_csr_pmp_7_cfg_a [0]}; 
    wire[31:0] core_csr_pmp_7_mask ={ core_csr_pmp_mask_base_7 [29:0]&~( core_csr_pmp_mask_base_7 [29:0]+30'h1),2'h3}; reg[31:0] core_csr_reg_misa ; 
    wire[1:0] core_csr_read_mstatus_lo_lo_lo_hi ={ core_csr_reg_mstatus_mie ,1'h0}; 
    wire[3:0] core_csr_read_mstatus_lo_lo_lo ={ core_csr_read_mstatus_lo_lo_lo_hi ,2'h0}; 
    wire[1:0] core_csr_read_mstatus_lo_lo_hi_hi_hi ={1'h0, core_csr_reg_mstatus_mpie }; 
    wire[2:0] core_csr_read_mstatus_lo_lo_hi_hi ={ core_csr_read_mstatus_lo_lo_hi_hi_hi ,1'h0}; 
    wire[4:0] core_csr_read_mstatus_lo_lo_hi ={ core_csr_read_mstatus_lo_lo_hi_hi ,2'h0}; 
    wire[8:0] core_csr_read_mstatus_lo_lo ={ core_csr_read_mstatus_lo_lo_hi , core_csr_read_mstatus_lo_lo_lo }; 
    wire[3:0] core_csr_read_mstatus_lo_hi_lo_lo ={ core_csr_reg_mstatus_mpp ,2'h0}; 
    wire[7:0] core_csr_read_mstatus_lo_hi_lo ={4'h0, core_csr_read_mstatus_lo_hi_lo_lo }; 
    wire[12:0] core_csr_read_mstatus_lo_hi ={5'h0, core_csr_read_mstatus_lo_hi_lo }; 
    wire[21:0] core_csr_read_mstatus_lo ={ core_csr_read_mstatus_lo_hi , core_csr_read_mstatus_lo_lo }; 
    wire[1:0] core_csr_read_mstatus_hi_lo_hi_hi_hi ={ core_csr_reg_mstatus_mpv , core_csr_reg_mstatus_gva }; 
    wire[2:0] core_csr_read_mstatus_hi_lo_hi_hi ={ core_csr_read_mstatus_hi_lo_hi_hi_hi ,1'h0}; 
    wire[5:0] core_csr_read_mstatus_hi_lo_hi ={ core_csr_read_mstatus_hi_lo_hi_hi ,3'h0}; 
    wire[17:0] core_csr_read_mstatus_hi_lo ={ core_csr_read_mstatus_hi_lo_hi ,12'h0}; 
    wire[2:0] core_csr_read_mstatus_hi_hi_lo_hi_hi ={ core_csr_reg_mstatus_v ,2'h3}; 
    wire[3:0] core_csr_read_mstatus_hi_hi_lo_hi ={ core_csr_read_mstatus_hi_hi_lo_hi_hi , core_csr_reg_mstatus_v }; 
    wire[27:0] core_csr_read_mstatus_hi_hi_lo ={ core_csr_read_mstatus_hi_hi_lo_hi ,24'h0}; 
    wire[33:0] core_csr_read_mstatus_hi_hi_hi_lo ={ core_csr_reg_misa ,2'h3}; 
    wire[1:0] core_csr_read_mstatus_hi_hi_hi_hi_hi ={ core_csr_reg_debug , core_csr_io_status_cease_r }; 
    wire[2:0] core_csr_read_mstatus_hi_hi_hi_hi ={ core_csr_read_mstatus_hi_hi_hi_hi_hi , core_csr_reg_wfi }; 
    wire[36:0] core_csr_read_mstatus_hi_hi_hi ={ core_csr_read_mstatus_hi_hi_hi_hi , core_csr_read_mstatus_hi_hi_hi_lo }; 
    wire[64:0] core_csr_read_mstatus_hi_hi ={ core_csr_read_mstatus_hi_hi_hi , core_csr_read_mstatus_hi_hi_lo }; 
    wire[82:0] core_csr_read_mstatus_hi ={ core_csr_read_mstatus_hi_hi , core_csr_read_mstatus_hi_lo }; 
    wire[31:0] core_csr_read_mstatus ={ core_csr_read_mstatus_hi [9:0], core_csr_read_mstatus_lo }; 
    wire[31:0] core_csr_read_mtvec = core_csr_reg_mtvec &{25'h1FFFFFF,~( core_csr_reg_mtvec [0] ? 7'h7E:7'h2)}; 
    wire[31:0] core_csr_notDebugTVec_base = core_csr_read_mtvec ; 
    wire[1:0] core_csr__GEN ={ core_csr_reg_bp_0_control_x , core_csr_reg_bp_0_control_w }; 
    wire[1:0] core_csr_lo_lo_hi_4 ; 
  assign  core_csr_lo_lo_hi_4 = core_csr__GEN ; 
    wire[1:0] core_csr_newBPC_lo_lo_hi ; 
  assign  core_csr_newBPC_lo_lo_hi = core_csr__GEN ; 
    wire[2:0] core_csr_lo_lo_4 ={ core_csr_lo_lo_hi_4 , core_csr_reg_bp_0_control_r }; 
    wire[6:0] core_csr_lo_4 ={4'h8, core_csr_lo_lo_4 }; 
    wire[3:0] core_csr__GEN_0 ={2'h0, core_csr_reg_bp_0_control_tmatch }; 
    wire[3:0] core_csr_hi_lo_lo_4 ; 
  assign  core_csr_hi_lo_lo_4 = core_csr__GEN_0 ; 
    wire[3:0] core_csr_newBPC_hi_lo_lo ; 
  assign  core_csr_newBPC_hi_lo_lo = core_csr__GEN_0 ; 
    wire[1:0] core_csr__GEN_1 ={ core_csr_reg_bp_0_control_action ,1'h0}; 
    wire[1:0] core_csr_hi_lo_hi_4 ; 
  assign  core_csr_hi_lo_hi_4 = core_csr__GEN_1 ; 
    wire[1:0] core_csr_newBPC_hi_lo_hi ; 
  assign  core_csr_newBPC_hi_lo_hi = core_csr__GEN_1 ; 
    wire[5:0] core_csr_hi_lo_4 ={ core_csr_hi_lo_hi_4 , core_csr_hi_lo_lo_4 }; 
    wire[4:0] core_csr__GEN_2 ={4'h2, core_csr_reg_bp_0_control_dmode }; 
    wire[4:0] core_csr_hi_hi_hi_4 ; 
  assign  core_csr_hi_hi_hi_4 = core_csr__GEN_2 ; 
    wire[4:0] core_csr_newBPC_hi_hi_hi ; 
  assign  core_csr_newBPC_hi_hi_hi = core_csr__GEN_2 ; 
    wire[18:0] core_csr_hi_hi_4 ={ core_csr_hi_hi_hi_4 ,14'h400}; 
    wire[24:0] core_csr_hi_4 ={ core_csr_hi_hi_4 , core_csr_hi_lo_4 }; 
    wire[1:0] core_csr_lo_5 ={ core_csr_lo_hi_5 ,1'h0}; 
    wire[31:0] core_csr__io_evec_T_20 =~ core_csr_reg_mepc ; 
    wire[1:0] core_csr__GEN_3 ={~( core_csr_reg_misa [2]),1'h1}; 
    wire[2:0] core_csr_lo_lo_hi_5 ={2'h0, core_csr_reg_dcsr_step }; 
    wire[4:0] core_csr_lo_lo_5 ={ core_csr_lo_lo_hi_5 ,2'h3}; 
    wire[3:0] core_csr_lo_hi_lo_5 ={ core_csr_reg_dcsr_cause , core_csr_reg_dcsr_v }; 
    wire[5:0] core_csr_lo_hi_6 ={2'h0, core_csr_lo_hi_lo_5 }; 
    wire[10:0] core_csr_lo_6 ={ core_csr_lo_hi_6 , core_csr_lo_lo_5 }; 
    wire[12:0] core_csr_hi_hi_lo_5 ={12'h0, core_csr_reg_dcsr_ebreakm }; 
    wire[16:0] core_csr_hi_hi_6 ={4'h4, core_csr_hi_hi_lo_5 }; 
    wire[20:0] core_csr_hi_6 ={ core_csr_hi_hi_6 ,4'h0}; 
    wire[31:0] core_csr__io_evec_T_10 =~ core_csr_reg_dpc ; 
    wire[1:0] core_csr_lo_hi_7 ={ core_csr_reg_pmp_0_cfg_x , core_csr_reg_pmp_0_cfg_w }; 
    wire[2:0] core_csr_lo_7 ={ core_csr_lo_hi_7 , core_csr_reg_pmp_0_cfg_r }; 
    wire[2:0] core_csr_hi_hi_7 ={ core_csr_reg_pmp_0_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_7 ={ core_csr_hi_hi_7 , core_csr_reg_pmp_0_cfg_a }; 
    wire[1:0] core_csr_lo_hi_8 ={ core_csr_reg_pmp_1_cfg_x , core_csr_reg_pmp_1_cfg_w }; 
    wire[2:0] core_csr_lo_8 ={ core_csr_lo_hi_8 , core_csr_reg_pmp_1_cfg_r }; 
    wire[2:0] core_csr_hi_hi_8 ={ core_csr_reg_pmp_1_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_8 ={ core_csr_hi_hi_8 , core_csr_reg_pmp_1_cfg_a }; 
    wire[1:0] core_csr_lo_hi_9 ={ core_csr_reg_pmp_2_cfg_x , core_csr_reg_pmp_2_cfg_w }; 
    wire[2:0] core_csr_lo_9 ={ core_csr_lo_hi_9 , core_csr_reg_pmp_2_cfg_r }; 
    wire[2:0] core_csr_hi_hi_9 ={ core_csr_reg_pmp_2_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_9 ={ core_csr_hi_hi_9 , core_csr_reg_pmp_2_cfg_a }; 
    wire[1:0] core_csr_lo_hi_10 ={ core_csr_reg_pmp_3_cfg_x , core_csr_reg_pmp_3_cfg_w }; 
    wire[2:0] core_csr_lo_10 ={ core_csr_lo_hi_10 , core_csr_reg_pmp_3_cfg_r }; 
    wire[2:0] core_csr_hi_hi_10 ={ core_csr_reg_pmp_3_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_10 ={ core_csr_hi_hi_10 , core_csr_reg_pmp_3_cfg_a }; 
    wire[15:0] core_csr_lo_11 ={ core_csr_hi_8 , core_csr_lo_8 , core_csr_hi_7 , core_csr_lo_7 }; 
    wire[15:0] core_csr_hi_11 ={ core_csr_hi_10 , core_csr_lo_10 , core_csr_hi_9 , core_csr_lo_9 }; 
    wire[1:0] core_csr_lo_hi_11 ={ core_csr_reg_pmp_4_cfg_x , core_csr_reg_pmp_4_cfg_w }; 
    wire[2:0] core_csr_lo_12 ={ core_csr_lo_hi_11 , core_csr_reg_pmp_4_cfg_r }; 
    wire[2:0] core_csr_hi_hi_11 ={ core_csr_reg_pmp_4_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_12 ={ core_csr_hi_hi_11 , core_csr_reg_pmp_4_cfg_a }; 
    wire[1:0] core_csr_lo_hi_12 ={ core_csr_reg_pmp_5_cfg_x , core_csr_reg_pmp_5_cfg_w }; 
    wire[2:0] core_csr_lo_13 ={ core_csr_lo_hi_12 , core_csr_reg_pmp_5_cfg_r }; 
    wire[2:0] core_csr_hi_hi_12 ={ core_csr_reg_pmp_5_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_13 ={ core_csr_hi_hi_12 , core_csr_reg_pmp_5_cfg_a }; 
    wire[1:0] core_csr_lo_hi_13 ={ core_csr_reg_pmp_6_cfg_x , core_csr_reg_pmp_6_cfg_w }; 
    wire[2:0] core_csr_lo_14 ={ core_csr_lo_hi_13 , core_csr_reg_pmp_6_cfg_r }; 
    wire[2:0] core_csr_hi_hi_13 ={ core_csr_reg_pmp_6_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_14 ={ core_csr_hi_hi_13 , core_csr_reg_pmp_6_cfg_a }; 
    wire[1:0] core_csr_lo_hi_14 ={ core_csr_reg_pmp_7_cfg_x , core_csr_reg_pmp_7_cfg_w }; 
    wire[2:0] core_csr_lo_15 ={ core_csr_lo_hi_14 , core_csr_reg_pmp_7_cfg_r }; 
    wire[2:0] core_csr_hi_hi_14 ={ core_csr_reg_pmp_7_cfg_l ,2'h0}; 
    wire[4:0] core_csr_hi_15 ={ core_csr_hi_hi_14 , core_csr_reg_pmp_7_cfg_a }; 
    wire[15:0] core_csr_lo_16 ={ core_csr_hi_13 , core_csr_lo_13 , core_csr_hi_12 , core_csr_lo_12 }; 
    wire[15:0] core_csr_hi_16 ={ core_csr_hi_15 , core_csr_lo_15 , core_csr_hi_14 , core_csr_lo_14 }; reg[31:0] core_csr_reg_custom_0 ; 
    wire core_csr_reg_custom_read =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'h7C1; 
    wire core_csr_reg_custom_read_1 =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'hF12; 
    wire core_csr_reg_custom_read_2 =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'hF11; 
    wire core_csr_reg_custom_read_3 =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'hF13; 
    wire[12:0] core_csr_addr ={ core_csr_reg_mstatus_v , core_csr_io_rw_addr }; 
    wire[11:0] core_csr_decoded_decoded_plaInput ; 
    wire[11:0] core_csr_decoded_decoded_invInputs =~ core_csr_decoded_decoded_plaInput ; 
    wire[195:0] core_csr_decoded_decoded_invMatrixOutputs ; 
    wire core_csr_decoded_decoded_andMatrixInput_0 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_2 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_6 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_8 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_10 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_12 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_14 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_16 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_18 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_20 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_22 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_24 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_26 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_28 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_30 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_32 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_34 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_36 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_39 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_41 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_43 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_45 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_47 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_49 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_51 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_53 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_55 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_57 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_59 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_61 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_63 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_68 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_70 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_72 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_74 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_76 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_78 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_80 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_82 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_84 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_86 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_88 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_90 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_92 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_94 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_96 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_99 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_101 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_103 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_105 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_107 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_109 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_111 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_113 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_115 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_117 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_119 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_121 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_123 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_125 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_127 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_130 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_132 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_134 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_136 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_138 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_140 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_142 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_144 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_146 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_148 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_150 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_152 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_154 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_156 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_158 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_161 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_163 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_165 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_167 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_169 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_171 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_173 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_175 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_177 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_179 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_181 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_183 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_185 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_187 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_189 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_192 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_194 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_1 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_2 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_3 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_4 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_6 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_7 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_10 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_11 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_14 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_15 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_18 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_19 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_22 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_23 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_26 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_27 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_30 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_31 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_34 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_35 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_39 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_40 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_43 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_44 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_47 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_48 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_51 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_52 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_55 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_56 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_59 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_60 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_63 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_64 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_67 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_70 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_71 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_74 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_75 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_78 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_79 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_82 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_83 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_86 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_87 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_90 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_91 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_94 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_95 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_98 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_101 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_102 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_105 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_106 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_109 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_110 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_113 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_114 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_117 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_118 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_121 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_122 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_125 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_126 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_129 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_132 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_133 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_136 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_137 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_140 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_141 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_144 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_145 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_148 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_149 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_152 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_153 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_156 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_157 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_160 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_163 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_164 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_167 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_168 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_171 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_172 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_175 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_176 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_179 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_180 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_183 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_184 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_187 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_188 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_191 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_194 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_195 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_1 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_4 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_5 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_10 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_11 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_12 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_13 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_18 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_19 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_20 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_21 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_26 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_27 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_28 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_29 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_34 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_35 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_36 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_37 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_39 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_40 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_41 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_42 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_43 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_44 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_45 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_46 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_51 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_52 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_53 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_54 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_59 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_60 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_61 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_62 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_63 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_64 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_65 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_67 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_68 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_69 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_74 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_75 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_76 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_77 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_82 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_83 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_84 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_85 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_90 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_91 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_92 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_93 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_98 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_99 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_100 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_105 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_106 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_107 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_108 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_113 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_114 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_115 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_116 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_121 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_122 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_123 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_124 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_129 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_130 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_131 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_136 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_137 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_138 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_139 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_144 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_145 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_146 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_147 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_152 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_153 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_154 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_155 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_160 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_161 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_162 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_167 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_168 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_169 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_170 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_175 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_176 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_177 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_178 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_183 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_184 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_185 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_186 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_191 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_192 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_193 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_1 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_2 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_3 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_4 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_5 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_6 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_7 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_8 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_9 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_18 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_19 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_20 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_21 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_22 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_23 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_24 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_25 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_34 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_35 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_36 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_37 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_38 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_39 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_40 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_41 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_42 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_43 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_44 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_45 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_46 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_47 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_48 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_49 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_50 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_59 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_60 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_61 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_62 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_63 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_64 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_65 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_67 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_68 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_69 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_70 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_71 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_72 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_73 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_82 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_83 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_84 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_85 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_86 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_87 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_88 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_89 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_98 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_99 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_100 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_101 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_102 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_103 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_104 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_113 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_114 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_115 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_116 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_117 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_118 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_119 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_120 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_129 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_130 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_131 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_132 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_133 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_134 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_135 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_144 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_145 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_146 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_147 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_148 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_149 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_150 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_151 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_160 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_161 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_162 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_163 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_164 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_165 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_166 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_175 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_176 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_177 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_178 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_179 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_180 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_181 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_182 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_191 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_192 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_193 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_194 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_195 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_1 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_2 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_3 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_4 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_5 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_6 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_7 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_8 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_9 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_10 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_11 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_12 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_13 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_14 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_15 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_16 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_17 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_34 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_35 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_36 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_37 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_38 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_39 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_40 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_41 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_42 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_59 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_60 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_61 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_62 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_67 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_68 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_69 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_70 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_71 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_72 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_73 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_74 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_75 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_76 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_77 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_78 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_79 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_80 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_81 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_98 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_99 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_100 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_101 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_102 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_103 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_104 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_105 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_106 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_107 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_108 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_109 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_110 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_111 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_112 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_129 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_130 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_131 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_132 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_133 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_134 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_135 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_136 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_137 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_138 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_139 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_140 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_141 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_142 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_143 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_160 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_161 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_162 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_163 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_164 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_165 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_166 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_167 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_168 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_169 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_170 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_171 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_172 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_173 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_174 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_1 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_2 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_3 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_34 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_35 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_36 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_37 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_38 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_67 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_68 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_69 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_70 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_71 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_72 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_73 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_74 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_75 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_76 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_77 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_78 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_79 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_80 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_81 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_82 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_83 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_84 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_85 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_86 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_87 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_88 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_89 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_90 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_91 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_92 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_93 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_94 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_95 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_96 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_97 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_98 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_99 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_100 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_101 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_102 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_103 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_104 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_105 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_106 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_107 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_108 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_109 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_110 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_111 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_112 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_113 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_114 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_115 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_116 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_117 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_118 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_119 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_120 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_121 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_122 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_123 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_124 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_125 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_126 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_127 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_128 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_129 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_130 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_131 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_132 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_133 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_134 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_135 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_136 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_137 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_138 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_139 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_140 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_141 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_142 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_143 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_144 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_145 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_146 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_147 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_148 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_149 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_150 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_151 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_152 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_153 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_154 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_155 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_156 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_157 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_158 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_159 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_160 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_161 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_162 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_163 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_164 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_165 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_166 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_167 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_168 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_169 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_170 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_171 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_172 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_173 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_174 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_175 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_176 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_177 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_178 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_179 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_180 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_181 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_182 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_183 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_184 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_185 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_186 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_187 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_188 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_189 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_190 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_191 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_192 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_193 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_194 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_195 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_1 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_2 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_3 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_4 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_5 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_6 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_7 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_8 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_9 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_10 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_11 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_12 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_13 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_14 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_15 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_16 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_17 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_18 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_19 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_20 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_21 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_22 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_23 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_24 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_25 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_26 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_27 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_28 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_29 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_30 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_31 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_32 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_33 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_39 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_40 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_41 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_42 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_43 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_44 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_45 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_46 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_47 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_48 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_49 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_50 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_51 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_52 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_53 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_54 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_55 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_56 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_57 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_58 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_59 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_60 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_61 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_62 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_63 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_64 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_65 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_67 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_67 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_68 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_69 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_70 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_71 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_72 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_73 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_74 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_75 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_76 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_77 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_78 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_79 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_80 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_81 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_82 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_83 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_84 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_85 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_86 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_87 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_88 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_89 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_90 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_91 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_92 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_93 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_94 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_95 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_96 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_98 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_98 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_99 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_100 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_101 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_102 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_103 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_104 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_105 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_106 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_107 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_108 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_109 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_110 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_111 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_112 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_113 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_114 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_115 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_116 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_117 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_118 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_119 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_120 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_121 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_122 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_123 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_124 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_125 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_126 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_127 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_129 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_129 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_130 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_131 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_132 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_133 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_134 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_135 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_136 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_137 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_138 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_139 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_140 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_141 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_142 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_143 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_144 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_145 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_146 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_147 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_148 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_149 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_150 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_151 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_152 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_153 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_154 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_155 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_156 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_157 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_158 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_160 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_160 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_161 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_162 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_163 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_164 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_165 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_166 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_167 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_168 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_169 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_170 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_171 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_172 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_173 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_174 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_175 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_176 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_177 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_178 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_179 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_180 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_181 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_182 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_183 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_184 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_185 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_186 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_187 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_188 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_189 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_191 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_191 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_192 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_193 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_194 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_1 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_2 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_3 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_4 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_5 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_6 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_7 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_8 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_9 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_10 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_11 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_12 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_13 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_14 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_15 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_16 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_17 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_18 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_19 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_20 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_21 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_22 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_23 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_24 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_25 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_26 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_27 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_28 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_29 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_30 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_31 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_32 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_33 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_34 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_35 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_36 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_37 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_38 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_66 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_67 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_68 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_69 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_70 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_71 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_72 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_73 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_74 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_75 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_76 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_77 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_78 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_79 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_80 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_81 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_82 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_83 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_84 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_85 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_86 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_87 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_88 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_89 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_90 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_91 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_92 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_93 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_94 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_95 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_96 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_128 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_129 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_130 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_131 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_132 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_133 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_134 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_135 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_136 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_137 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_138 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_139 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_140 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_141 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_142 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_143 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_144 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_145 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_146 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_147 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_148 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_149 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_150 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_151 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_152 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_153 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_154 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_155 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_156 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_157 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_158 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_190 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_191 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_192 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_193 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_194 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_1 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_2 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_3 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_4 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_5 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_6 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_7 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_8 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_9 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_10 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_11 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_12 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_13 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_14 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_15 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_16 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_17 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_18 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_19 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_20 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_21 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_22 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_23 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_24 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_25 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_26 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_27 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_28 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_29 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_30 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_31 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_32 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_33 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_34 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_35 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_36 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_37 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_38 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_39 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_40 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_41 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_42 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_43 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_44 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_45 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_46 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_47 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_48 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_49 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_50 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_51 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_52 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_53 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_54 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_55 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_56 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_57 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_58 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_59 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_60 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_61 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_62 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_63 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_64 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_65 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_66 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_66 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_67 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_68 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_69 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_70 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_71 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_72 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_73 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_74 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_75 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_76 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_77 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_78 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_79 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_80 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_81 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_82 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_83 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_84 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_85 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_86 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_87 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_88 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_89 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_90 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_91 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_92 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_93 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_94 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_95 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_96 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_97 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_98 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_99 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_100 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_101 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_102 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_103 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_104 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_105 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_106 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_107 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_108 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_109 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_110 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_111 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_112 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_113 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_114 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_115 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_116 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_117 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_118 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_119 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_120 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_121 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_122 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_123 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_124 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_125 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_126 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_127 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_190 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_191 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_192 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_193 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_194 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_1 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_2 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_3 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_4 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_5 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_6 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_7 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_8 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_9 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_10 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_11 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_12 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_13 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_14 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_15 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_16 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_17 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_18 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_19 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_20 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_21 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_22 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_23 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_24 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_25 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_26 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_27 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_28 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_29 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_30 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_31 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_32 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_33 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_34 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_35 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_36 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_37 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_38 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_39 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_40 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_41 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_42 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_43 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_44 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_45 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_46 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_47 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_48 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_49 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_50 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_51 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_52 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_53 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_54 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_55 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_56 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_57 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_58 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_59 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_60 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_61 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_62 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_63 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_64 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_65 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_66 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_66 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_67 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_68 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_69 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_70 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_71 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_72 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_73 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_74 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_75 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_76 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_77 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_78 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_79 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_80 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_81 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_82 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_83 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_84 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_85 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_86 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_87 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_88 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_89 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_90 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_91 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_92 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_93 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_94 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_95 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_96 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_97 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_98 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_99 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_100 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_101 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_102 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_103 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_104 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_105 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_106 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_107 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_108 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_109 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_110 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_111 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_112 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_113 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_114 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_115 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_116 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_117 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_118 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_119 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_120 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_121 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_122 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_123 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_124 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_125 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_126 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_127 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_190 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_191 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_192 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_193 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_194 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_1 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_2 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_3 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_4 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_5 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_6 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_7 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_8 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_9 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_10 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_11 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_12 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_13 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_14 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_15 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_16 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_17 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_18 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_19 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_20 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_21 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_22 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_23 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_24 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_25 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_26 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_27 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_28 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_29 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_30 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_31 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_32 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_33 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_34 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_35 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_36 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_37 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_38 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_38 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_39 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_40 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_41 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_42 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_43 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_44 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_45 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_46 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_47 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_48 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_49 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_50 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_51 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_52 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_53 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_54 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_55 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_56 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_57 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_66 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_66 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_67 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_68 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_69 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_70 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_71 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_72 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_73 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_74 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_75 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_76 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_77 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_78 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_79 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_80 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_81 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_82 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_83 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_84 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_85 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_86 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_87 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_88 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_89 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_90 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_91 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_92 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_93 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_94 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_95 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_97 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_97 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_98 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_99 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_100 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_101 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_102 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_103 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_104 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_105 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_106 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_107 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_108 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_109 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_110 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_111 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_112 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_113 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_114 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_115 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_116 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_117 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_118 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_119 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_120 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_121 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_122 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_123 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_124 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_125 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_126 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_1 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_2 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_3 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_4 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_5 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_4 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_5 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_6 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_7 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_8 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_9 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_10 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_11 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_12 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_13 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_14 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_15 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_16 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_17 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_18 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_19 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_20 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_21 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_22 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_23 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_24 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_25 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_26 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_27 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_28 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_29 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_30 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_31 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_32 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_33 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_34 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_35 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_38 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_36 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_37 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_38 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_39 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_40 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_41 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_42 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_43 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_44 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_45 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_46 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_47 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_48 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_49 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_50 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_51 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_52 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_53 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_54 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_55 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_56 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_57 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_58 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_59 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_60 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_61 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_64 = core_csr_decoded_decoded_invInputs [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_66 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi ={ core_csr_decoded_decoded_andMatrixInput_9 , core_csr_decoded_decoded_andMatrixInput_10 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo ={ core_csr_decoded_decoded_lo_lo_hi , core_csr_decoded_decoded_andMatrixInput_11 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi ={ core_csr_decoded_decoded_andMatrixInput_6 , core_csr_decoded_decoded_andMatrixInput_7 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi ={ core_csr_decoded_decoded_lo_hi_hi , core_csr_decoded_decoded_andMatrixInput_8 }; 
    wire[5:0] core_csr_decoded_decoded_lo ={ core_csr_decoded_decoded_lo_hi , core_csr_decoded_decoded_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi ={ core_csr_decoded_decoded_andMatrixInput_3 , core_csr_decoded_decoded_andMatrixInput_4 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo ={ core_csr_decoded_decoded_hi_lo_hi , core_csr_decoded_decoded_andMatrixInput_5 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi ={ core_csr_decoded_decoded_andMatrixInput_0 , core_csr_decoded_decoded_andMatrixInput_1 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi ={ core_csr_decoded_decoded_hi_hi_hi , core_csr_decoded_decoded_andMatrixInput_2 }; 
    wire[5:0] core_csr_decoded_decoded_hi ={ core_csr_decoded_decoded_hi_hi , core_csr_decoded_decoded_hi_lo }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_1 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_3 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_7 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_9 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_11 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_13 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_15 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_17 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_19 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_21 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_23 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_25 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_27 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_29 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_31 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_33 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_35 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_37 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_40 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_42 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_44 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_46 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_48 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_50 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_52 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_54 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_56 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_58 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_60 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_62 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_64 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_69 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_71 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_73 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_75 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_77 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_79 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_81 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_83 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_85 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_87 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_89 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_91 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_93 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_95 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_97 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_100 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_102 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_104 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_106 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_108 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_110 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_112 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_114 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_116 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_118 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_120 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_122 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_124 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_126 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_128 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_131 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_133 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_135 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_137 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_139 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_141 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_143 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_145 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_147 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_149 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_151 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_153 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_155 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_157 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_159 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_162 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_164 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_166 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_168 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_170 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_172 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_174 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_176 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_178 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_180 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_182 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_184 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_186 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_188 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_190 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_193 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_195 = core_csr_decoded_decoded_plaInput [0]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_9_1 , core_csr_decoded_decoded_andMatrixInput_10_1 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_1 ={ core_csr_decoded_decoded_lo_lo_hi_1 , core_csr_decoded_decoded_andMatrixInput_11_1 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_6_1 , core_csr_decoded_decoded_andMatrixInput_7_1 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_1 ={ core_csr_decoded_decoded_lo_hi_hi_1 , core_csr_decoded_decoded_andMatrixInput_8_1 }; 
    wire[5:0] core_csr_decoded_decoded_lo_1 ={ core_csr_decoded_decoded_lo_hi_1 , core_csr_decoded_decoded_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_3_1 , core_csr_decoded_decoded_andMatrixInput_4_1 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_1 ={ core_csr_decoded_decoded_hi_lo_hi_1 , core_csr_decoded_decoded_andMatrixInput_5_1 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_0_1 , core_csr_decoded_decoded_andMatrixInput_1_1 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_1 ={ core_csr_decoded_decoded_hi_hi_hi_1 , core_csr_decoded_decoded_andMatrixInput_2_1 }; 
    wire[5:0] core_csr_decoded_decoded_hi_1 ={ core_csr_decoded_decoded_hi_hi_1 , core_csr_decoded_decoded_hi_lo_1 }; 
    wire core_csr_decoded_decoded_andMatrixInput_2_2 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_3 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_6 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_7 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_8 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_9 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_14 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_15 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_16 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_17 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_22 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_23 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_24 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_25 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_30 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_31 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_32 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_33 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_38 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_47 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_48 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_49 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_50 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_55 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_56 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_57 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_58 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_70 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_71 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_72 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_73 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_78 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_79 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_80 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_81 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_86 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_87 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_88 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_89 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_94 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_95 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_96 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_97 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_101 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_102 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_103 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_104 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_109 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_110 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_111 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_112 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_117 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_118 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_119 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_120 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_125 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_126 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_127 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_128 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_132 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_133 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_134 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_135 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_140 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_141 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_142 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_143 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_148 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_149 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_150 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_151 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_156 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_157 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_158 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_159 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_163 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_164 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_165 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_166 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_171 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_172 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_173 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_174 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_179 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_180 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_181 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_182 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_187 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_188 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_189 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_190 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_194 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_195 = core_csr_decoded_decoded_plaInput [2]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_9_2 , core_csr_decoded_decoded_andMatrixInput_10_2 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_2 ={ core_csr_decoded_decoded_lo_lo_hi_2 , core_csr_decoded_decoded_andMatrixInput_11_2 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_6_2 , core_csr_decoded_decoded_andMatrixInput_7_2 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_2 ={ core_csr_decoded_decoded_lo_hi_hi_2 , core_csr_decoded_decoded_andMatrixInput_8_2 }; 
    wire[5:0] core_csr_decoded_decoded_lo_2 ={ core_csr_decoded_decoded_lo_hi_2 , core_csr_decoded_decoded_lo_lo_2 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_3_2 , core_csr_decoded_decoded_andMatrixInput_4_2 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_2 ={ core_csr_decoded_decoded_hi_lo_hi_2 , core_csr_decoded_decoded_andMatrixInput_5_2 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_0_2 , core_csr_decoded_decoded_andMatrixInput_1_2 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_2 ={ core_csr_decoded_decoded_hi_hi_hi_2 , core_csr_decoded_decoded_andMatrixInput_2_2 }; 
    wire[5:0] core_csr_decoded_decoded_hi_2 ={ core_csr_decoded_decoded_hi_hi_2 , core_csr_decoded_decoded_hi_lo_2 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_9_3 , core_csr_decoded_decoded_andMatrixInput_10_3 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_3 ={ core_csr_decoded_decoded_lo_lo_hi_3 , core_csr_decoded_decoded_andMatrixInput_11_3 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_6_3 , core_csr_decoded_decoded_andMatrixInput_7_3 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_3 ={ core_csr_decoded_decoded_lo_hi_hi_3 , core_csr_decoded_decoded_andMatrixInput_8_3 }; 
    wire[5:0] core_csr_decoded_decoded_lo_3 ={ core_csr_decoded_decoded_lo_hi_3 , core_csr_decoded_decoded_lo_lo_3 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_3_3 , core_csr_decoded_decoded_andMatrixInput_4_3 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_3 ={ core_csr_decoded_decoded_hi_lo_hi_3 , core_csr_decoded_decoded_andMatrixInput_5_3 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_0_3 , core_csr_decoded_decoded_andMatrixInput_1_3 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_3 ={ core_csr_decoded_decoded_hi_hi_hi_3 , core_csr_decoded_decoded_andMatrixInput_2_3 }; 
    wire[5:0] core_csr_decoded_decoded_hi_3 ={ core_csr_decoded_decoded_hi_hi_3 , core_csr_decoded_decoded_hi_lo_3 }; 
    wire core_csr_decoded_decoded_andMatrixInput_4_4 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_5 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_6 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_7 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_8 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_9 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_10 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_11 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_12 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_13 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_14 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_15 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_16 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_17 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_18 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_19 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_20 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_21 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_22 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_23 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_24 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_25 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_26 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_27 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_28 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_29 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_30 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_31 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_32 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_33 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_39 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_40 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_41 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_42 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_43 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_44 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_45 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_46 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_47 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_48 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_49 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_50 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_51 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_52 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_53 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_54 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_55 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_56 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_57 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_58 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_59 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_60 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_61 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_62 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_63 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_64 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_65 = core_csr_decoded_decoded_plaInput [5]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_4 ={ core_csr_decoded_decoded_andMatrixInput_9_4 , core_csr_decoded_decoded_andMatrixInput_10_4 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_6_4 , core_csr_decoded_decoded_andMatrixInput_7_4 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_4 ={ core_csr_decoded_decoded_lo_hi_hi_4 , core_csr_decoded_decoded_andMatrixInput_8_4 }; 
    wire[4:0] core_csr_decoded_decoded_lo_4 ={ core_csr_decoded_decoded_lo_hi_4 , core_csr_decoded_decoded_lo_lo_4 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_3_4 , core_csr_decoded_decoded_andMatrixInput_4_4 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_4 ={ core_csr_decoded_decoded_hi_lo_hi_4 , core_csr_decoded_decoded_andMatrixInput_5_4 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_0_4 , core_csr_decoded_decoded_andMatrixInput_1_4 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_4 ={ core_csr_decoded_decoded_hi_hi_hi_4 , core_csr_decoded_decoded_andMatrixInput_2_4 }; 
    wire[5:0] core_csr_decoded_decoded_hi_4 ={ core_csr_decoded_decoded_hi_hi_4 , core_csr_decoded_decoded_hi_lo_4 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_5 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_8 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_9 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_12 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_13 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_16 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_17 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_20 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_21 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_24 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_25 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_28 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_29 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_32 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_33 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_36 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_37 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_41 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_42 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_45 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_46 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_49 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_50 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_53 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_54 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_57 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_58 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_61 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_62 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_65 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_68 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_69 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_72 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_73 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_76 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_77 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_80 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_81 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_84 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_85 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_88 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_89 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_92 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_93 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_96 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_97 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_99 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_100 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_103 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_104 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_107 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_108 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_111 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_112 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_115 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_116 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_119 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_120 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_123 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_124 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_127 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_128 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_130 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_131 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_134 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_135 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_138 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_139 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_142 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_143 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_146 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_147 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_150 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_151 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_154 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_155 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_158 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_159 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_161 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_162 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_165 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_166 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_169 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_170 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_173 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_174 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_177 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_178 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_181 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_182 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_185 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_186 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_189 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_190 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_192 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_193 = core_csr_decoded_decoded_plaInput [1]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_5 ={ core_csr_decoded_decoded_andMatrixInput_9_5 , core_csr_decoded_decoded_andMatrixInput_10_5 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_6_5 , core_csr_decoded_decoded_andMatrixInput_7_5 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_5 ={ core_csr_decoded_decoded_lo_hi_hi_5 , core_csr_decoded_decoded_andMatrixInput_8_5 }; 
    wire[4:0] core_csr_decoded_decoded_lo_5 ={ core_csr_decoded_decoded_lo_hi_5 , core_csr_decoded_decoded_lo_lo_5 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_3_5 , core_csr_decoded_decoded_andMatrixInput_4_5 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_5 ={ core_csr_decoded_decoded_hi_lo_hi_5 , core_csr_decoded_decoded_andMatrixInput_5_5 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_0_5 , core_csr_decoded_decoded_andMatrixInput_1_5 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_5 ={ core_csr_decoded_decoded_hi_hi_hi_5 , core_csr_decoded_decoded_andMatrixInput_2_5 }; 
    wire[5:0] core_csr_decoded_decoded_hi_5 ={ core_csr_decoded_decoded_hi_hi_5 , core_csr_decoded_decoded_hi_lo_5 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_9_6 , core_csr_decoded_decoded_andMatrixInput_10_6 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_6 ={ core_csr_decoded_decoded_lo_lo_hi_4 , core_csr_decoded_decoded_andMatrixInput_11_4 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_6_6 , core_csr_decoded_decoded_andMatrixInput_7_6 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_6 ={ core_csr_decoded_decoded_lo_hi_hi_6 , core_csr_decoded_decoded_andMatrixInput_8_6 }; 
    wire[5:0] core_csr_decoded_decoded_lo_6 ={ core_csr_decoded_decoded_lo_hi_6 , core_csr_decoded_decoded_lo_lo_6 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_3_6 , core_csr_decoded_decoded_andMatrixInput_4_6 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_6 ={ core_csr_decoded_decoded_hi_lo_hi_6 , core_csr_decoded_decoded_andMatrixInput_5_6 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_0_6 , core_csr_decoded_decoded_andMatrixInput_1_6 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_6 ={ core_csr_decoded_decoded_hi_hi_hi_6 , core_csr_decoded_decoded_andMatrixInput_2_6 }; 
    wire[5:0] core_csr_decoded_decoded_hi_6 ={ core_csr_decoded_decoded_hi_hi_6 , core_csr_decoded_decoded_hi_lo_6 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_9_7 , core_csr_decoded_decoded_andMatrixInput_10_7 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_7 ={ core_csr_decoded_decoded_lo_lo_hi_5 , core_csr_decoded_decoded_andMatrixInput_11_5 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_6_7 , core_csr_decoded_decoded_andMatrixInput_7_7 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_7 ={ core_csr_decoded_decoded_lo_hi_hi_7 , core_csr_decoded_decoded_andMatrixInput_8_7 }; 
    wire[5:0] core_csr_decoded_decoded_lo_7 ={ core_csr_decoded_decoded_lo_hi_7 , core_csr_decoded_decoded_lo_lo_7 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_3_7 , core_csr_decoded_decoded_andMatrixInput_4_7 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_7 ={ core_csr_decoded_decoded_hi_lo_hi_7 , core_csr_decoded_decoded_andMatrixInput_5_7 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_0_7 , core_csr_decoded_decoded_andMatrixInput_1_7 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_7 ={ core_csr_decoded_decoded_hi_hi_hi_7 , core_csr_decoded_decoded_andMatrixInput_2_7 }; 
    wire[5:0] core_csr_decoded_decoded_hi_7 ={ core_csr_decoded_decoded_hi_hi_7 , core_csr_decoded_decoded_hi_lo_7 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_9_8 , core_csr_decoded_decoded_andMatrixInput_10_8 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_8 ={ core_csr_decoded_decoded_lo_lo_hi_6 , core_csr_decoded_decoded_andMatrixInput_11_6 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_6_8 , core_csr_decoded_decoded_andMatrixInput_7_8 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_8 ={ core_csr_decoded_decoded_lo_hi_hi_8 , core_csr_decoded_decoded_andMatrixInput_8_8 }; 
    wire[5:0] core_csr_decoded_decoded_lo_8 ={ core_csr_decoded_decoded_lo_hi_8 , core_csr_decoded_decoded_lo_lo_8 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_3_8 , core_csr_decoded_decoded_andMatrixInput_4_8 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_8 ={ core_csr_decoded_decoded_hi_lo_hi_8 , core_csr_decoded_decoded_andMatrixInput_5_8 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_0_8 , core_csr_decoded_decoded_andMatrixInput_1_8 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_8 ={ core_csr_decoded_decoded_hi_hi_hi_8 , core_csr_decoded_decoded_andMatrixInput_2_8 }; 
    wire[5:0] core_csr_decoded_decoded_hi_8 ={ core_csr_decoded_decoded_hi_hi_8 , core_csr_decoded_decoded_hi_lo_8 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_9_9 , core_csr_decoded_decoded_andMatrixInput_10_9 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_9 ={ core_csr_decoded_decoded_lo_lo_hi_7 , core_csr_decoded_decoded_andMatrixInput_11_7 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_6_9 , core_csr_decoded_decoded_andMatrixInput_7_9 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_9 ={ core_csr_decoded_decoded_lo_hi_hi_9 , core_csr_decoded_decoded_andMatrixInput_8_9 }; 
    wire[5:0] core_csr_decoded_decoded_lo_9 ={ core_csr_decoded_decoded_lo_hi_9 , core_csr_decoded_decoded_lo_lo_9 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_3_9 , core_csr_decoded_decoded_andMatrixInput_4_9 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_9 ={ core_csr_decoded_decoded_hi_lo_hi_9 , core_csr_decoded_decoded_andMatrixInput_5_9 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_0_9 , core_csr_decoded_decoded_andMatrixInput_1_9 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_9 ={ core_csr_decoded_decoded_hi_hi_hi_9 , core_csr_decoded_decoded_andMatrixInput_2_9 }; 
    wire[5:0] core_csr_decoded_decoded_hi_9 ={ core_csr_decoded_decoded_hi_hi_9 , core_csr_decoded_decoded_hi_lo_9 }; 
    wire core_csr_decoded_decoded_andMatrixInput_3_10 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_11 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_12 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_13 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_14 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_15 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_16 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_17 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_26 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_27 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_28 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_29 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_30 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_31 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_32 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_33 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_51 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_52 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_53 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_54 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_55 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_56 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_57 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_58 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_74 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_75 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_76 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_77 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_78 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_79 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_80 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_81 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_90 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_91 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_92 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_93 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_94 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_95 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_96 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_97 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_105 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_106 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_107 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_108 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_109 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_110 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_111 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_112 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_121 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_122 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_123 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_124 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_125 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_126 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_127 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_128 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_136 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_137 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_138 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_139 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_140 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_141 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_142 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_143 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_152 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_153 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_154 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_155 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_156 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_157 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_158 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_159 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_167 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_168 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_169 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_170 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_171 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_172 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_173 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_174 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_183 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_184 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_185 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_186 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_187 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_188 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_189 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_190 = core_csr_decoded_decoded_plaInput [3]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_9_10 , core_csr_decoded_decoded_andMatrixInput_10_10 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_10 ={ core_csr_decoded_decoded_lo_lo_hi_8 , core_csr_decoded_decoded_andMatrixInput_11_8 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_6_10 , core_csr_decoded_decoded_andMatrixInput_7_10 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_10 ={ core_csr_decoded_decoded_lo_hi_hi_10 , core_csr_decoded_decoded_andMatrixInput_8_10 }; 
    wire[5:0] core_csr_decoded_decoded_lo_10 ={ core_csr_decoded_decoded_lo_hi_10 , core_csr_decoded_decoded_lo_lo_10 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_3_10 , core_csr_decoded_decoded_andMatrixInput_4_10 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_10 ={ core_csr_decoded_decoded_hi_lo_hi_10 , core_csr_decoded_decoded_andMatrixInput_5_10 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_0_10 , core_csr_decoded_decoded_andMatrixInput_1_10 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_10 ={ core_csr_decoded_decoded_hi_hi_hi_10 , core_csr_decoded_decoded_andMatrixInput_2_10 }; 
    wire[5:0] core_csr_decoded_decoded_hi_10 ={ core_csr_decoded_decoded_hi_hi_10 , core_csr_decoded_decoded_hi_lo_10 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_9_11 , core_csr_decoded_decoded_andMatrixInput_10_11 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_11 ={ core_csr_decoded_decoded_lo_lo_hi_9 , core_csr_decoded_decoded_andMatrixInput_11_9 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_6_11 , core_csr_decoded_decoded_andMatrixInput_7_11 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_11 ={ core_csr_decoded_decoded_lo_hi_hi_11 , core_csr_decoded_decoded_andMatrixInput_8_11 }; 
    wire[5:0] core_csr_decoded_decoded_lo_11 ={ core_csr_decoded_decoded_lo_hi_11 , core_csr_decoded_decoded_lo_lo_11 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_3_11 , core_csr_decoded_decoded_andMatrixInput_4_11 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_11 ={ core_csr_decoded_decoded_hi_lo_hi_11 , core_csr_decoded_decoded_andMatrixInput_5_11 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_0_11 , core_csr_decoded_decoded_andMatrixInput_1_11 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_11 ={ core_csr_decoded_decoded_hi_hi_hi_11 , core_csr_decoded_decoded_andMatrixInput_2_11 }; 
    wire[5:0] core_csr_decoded_decoded_hi_11 ={ core_csr_decoded_decoded_hi_hi_11 , core_csr_decoded_decoded_hi_lo_11 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_9_12 , core_csr_decoded_decoded_andMatrixInput_10_12 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_12 ={ core_csr_decoded_decoded_lo_lo_hi_10 , core_csr_decoded_decoded_andMatrixInput_11_10 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_6_12 , core_csr_decoded_decoded_andMatrixInput_7_12 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_12 ={ core_csr_decoded_decoded_lo_hi_hi_12 , core_csr_decoded_decoded_andMatrixInput_8_12 }; 
    wire[5:0] core_csr_decoded_decoded_lo_12 ={ core_csr_decoded_decoded_lo_hi_12 , core_csr_decoded_decoded_lo_lo_12 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_3_12 , core_csr_decoded_decoded_andMatrixInput_4_12 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_12 ={ core_csr_decoded_decoded_hi_lo_hi_12 , core_csr_decoded_decoded_andMatrixInput_5_12 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_0_12 , core_csr_decoded_decoded_andMatrixInput_1_12 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_12 ={ core_csr_decoded_decoded_hi_hi_hi_12 , core_csr_decoded_decoded_andMatrixInput_2_12 }; 
    wire[5:0] core_csr_decoded_decoded_hi_12 ={ core_csr_decoded_decoded_hi_hi_12 , core_csr_decoded_decoded_hi_lo_12 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_9_13 , core_csr_decoded_decoded_andMatrixInput_10_13 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_13 ={ core_csr_decoded_decoded_lo_lo_hi_11 , core_csr_decoded_decoded_andMatrixInput_11_11 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_6_13 , core_csr_decoded_decoded_andMatrixInput_7_13 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_13 ={ core_csr_decoded_decoded_lo_hi_hi_13 , core_csr_decoded_decoded_andMatrixInput_8_13 }; 
    wire[5:0] core_csr_decoded_decoded_lo_13 ={ core_csr_decoded_decoded_lo_hi_13 , core_csr_decoded_decoded_lo_lo_13 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_3_13 , core_csr_decoded_decoded_andMatrixInput_4_13 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_13 ={ core_csr_decoded_decoded_hi_lo_hi_13 , core_csr_decoded_decoded_andMatrixInput_5_13 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_0_13 , core_csr_decoded_decoded_andMatrixInput_1_13 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_13 ={ core_csr_decoded_decoded_hi_hi_hi_13 , core_csr_decoded_decoded_andMatrixInput_2_13 }; 
    wire[5:0] core_csr_decoded_decoded_hi_13 ={ core_csr_decoded_decoded_hi_hi_13 , core_csr_decoded_decoded_hi_lo_13 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_9_14 , core_csr_decoded_decoded_andMatrixInput_10_14 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_14 ={ core_csr_decoded_decoded_lo_lo_hi_12 , core_csr_decoded_decoded_andMatrixInput_11_12 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_6_14 , core_csr_decoded_decoded_andMatrixInput_7_14 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_14 ={ core_csr_decoded_decoded_lo_hi_hi_14 , core_csr_decoded_decoded_andMatrixInput_8_14 }; 
    wire[5:0] core_csr_decoded_decoded_lo_14 ={ core_csr_decoded_decoded_lo_hi_14 , core_csr_decoded_decoded_lo_lo_14 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_3_14 , core_csr_decoded_decoded_andMatrixInput_4_14 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_14 ={ core_csr_decoded_decoded_hi_lo_hi_14 , core_csr_decoded_decoded_andMatrixInput_5_14 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_0_14 , core_csr_decoded_decoded_andMatrixInput_1_14 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_14 ={ core_csr_decoded_decoded_hi_hi_hi_14 , core_csr_decoded_decoded_andMatrixInput_2_14 }; 
    wire[5:0] core_csr_decoded_decoded_hi_14 ={ core_csr_decoded_decoded_hi_hi_14 , core_csr_decoded_decoded_hi_lo_14 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_9_15 , core_csr_decoded_decoded_andMatrixInput_10_15 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_15 ={ core_csr_decoded_decoded_lo_lo_hi_13 , core_csr_decoded_decoded_andMatrixInput_11_13 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_6_15 , core_csr_decoded_decoded_andMatrixInput_7_15 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_15 ={ core_csr_decoded_decoded_lo_hi_hi_15 , core_csr_decoded_decoded_andMatrixInput_8_15 }; 
    wire[5:0] core_csr_decoded_decoded_lo_15 ={ core_csr_decoded_decoded_lo_hi_15 , core_csr_decoded_decoded_lo_lo_15 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_3_15 , core_csr_decoded_decoded_andMatrixInput_4_15 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_15 ={ core_csr_decoded_decoded_hi_lo_hi_15 , core_csr_decoded_decoded_andMatrixInput_5_15 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_0_15 , core_csr_decoded_decoded_andMatrixInput_1_15 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_15 ={ core_csr_decoded_decoded_hi_hi_hi_15 , core_csr_decoded_decoded_andMatrixInput_2_15 }; 
    wire[5:0] core_csr_decoded_decoded_hi_15 ={ core_csr_decoded_decoded_hi_hi_15 , core_csr_decoded_decoded_hi_lo_15 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_9_16 , core_csr_decoded_decoded_andMatrixInput_10_16 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_16 ={ core_csr_decoded_decoded_lo_lo_hi_14 , core_csr_decoded_decoded_andMatrixInput_11_14 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_6_16 , core_csr_decoded_decoded_andMatrixInput_7_16 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_16 ={ core_csr_decoded_decoded_lo_hi_hi_16 , core_csr_decoded_decoded_andMatrixInput_8_16 }; 
    wire[5:0] core_csr_decoded_decoded_lo_16 ={ core_csr_decoded_decoded_lo_hi_16 , core_csr_decoded_decoded_lo_lo_16 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_3_16 , core_csr_decoded_decoded_andMatrixInput_4_16 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_16 ={ core_csr_decoded_decoded_hi_lo_hi_16 , core_csr_decoded_decoded_andMatrixInput_5_16 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_0_16 , core_csr_decoded_decoded_andMatrixInput_1_16 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_16 ={ core_csr_decoded_decoded_hi_hi_hi_16 , core_csr_decoded_decoded_andMatrixInput_2_16 }; 
    wire[5:0] core_csr_decoded_decoded_hi_16 ={ core_csr_decoded_decoded_hi_hi_16 , core_csr_decoded_decoded_hi_lo_16 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_9_17 , core_csr_decoded_decoded_andMatrixInput_10_17 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_17 ={ core_csr_decoded_decoded_lo_lo_hi_15 , core_csr_decoded_decoded_andMatrixInput_11_15 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_6_17 , core_csr_decoded_decoded_andMatrixInput_7_17 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_17 ={ core_csr_decoded_decoded_lo_hi_hi_17 , core_csr_decoded_decoded_andMatrixInput_8_17 }; 
    wire[5:0] core_csr_decoded_decoded_lo_17 ={ core_csr_decoded_decoded_lo_hi_17 , core_csr_decoded_decoded_lo_lo_17 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_3_17 , core_csr_decoded_decoded_andMatrixInput_4_17 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_17 ={ core_csr_decoded_decoded_hi_lo_hi_17 , core_csr_decoded_decoded_andMatrixInput_5_17 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_0_17 , core_csr_decoded_decoded_andMatrixInput_1_17 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_17 ={ core_csr_decoded_decoded_hi_hi_hi_17 , core_csr_decoded_decoded_andMatrixInput_2_17 }; 
    wire[5:0] core_csr_decoded_decoded_hi_17 ={ core_csr_decoded_decoded_hi_hi_17 , core_csr_decoded_decoded_hi_lo_17 }; 
    wire core_csr_decoded_decoded_andMatrixInput_4_18 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_19 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_20 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_21 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_22 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_23 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_24 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_25 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_26 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_27 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_28 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_29 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_30 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_31 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_32 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_33 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_43 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_44 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_45 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_46 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_47 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_48 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_49 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_50 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_51 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_52 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_53 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_54 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_55 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_56 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_57 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_58 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_63 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_64 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_65 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_82 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_83 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_84 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_85 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_86 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_87 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_88 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_89 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_90 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_91 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_92 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_93 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_94 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_95 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_96 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_97 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_113 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_114 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_115 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_116 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_117 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_118 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_119 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_120 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_121 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_122 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_123 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_124 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_125 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_126 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_127 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_128 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_144 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_145 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_146 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_147 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_148 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_149 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_150 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_151 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_152 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_153 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_154 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_155 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_156 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_157 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_158 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_159 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_175 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_176 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_177 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_178 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_179 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_180 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_181 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_182 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_183 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_184 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_185 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_186 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_187 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_188 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_189 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_190 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_191 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_192 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_193 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_194 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_195 = core_csr_decoded_decoded_plaInput [4]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_9_18 , core_csr_decoded_decoded_andMatrixInput_10_18 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_18 ={ core_csr_decoded_decoded_lo_lo_hi_16 , core_csr_decoded_decoded_andMatrixInput_11_16 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_6_18 , core_csr_decoded_decoded_andMatrixInput_7_18 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_18 ={ core_csr_decoded_decoded_lo_hi_hi_18 , core_csr_decoded_decoded_andMatrixInput_8_18 }; 
    wire[5:0] core_csr_decoded_decoded_lo_18 ={ core_csr_decoded_decoded_lo_hi_18 , core_csr_decoded_decoded_lo_lo_18 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_3_18 , core_csr_decoded_decoded_andMatrixInput_4_18 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_18 ={ core_csr_decoded_decoded_hi_lo_hi_18 , core_csr_decoded_decoded_andMatrixInput_5_18 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_0_18 , core_csr_decoded_decoded_andMatrixInput_1_18 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_18 ={ core_csr_decoded_decoded_hi_hi_hi_18 , core_csr_decoded_decoded_andMatrixInput_2_18 }; 
    wire[5:0] core_csr_decoded_decoded_hi_18 ={ core_csr_decoded_decoded_hi_hi_18 , core_csr_decoded_decoded_hi_lo_18 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_9_19 , core_csr_decoded_decoded_andMatrixInput_10_19 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_19 ={ core_csr_decoded_decoded_lo_lo_hi_17 , core_csr_decoded_decoded_andMatrixInput_11_17 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_6_19 , core_csr_decoded_decoded_andMatrixInput_7_19 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_19 ={ core_csr_decoded_decoded_lo_hi_hi_19 , core_csr_decoded_decoded_andMatrixInput_8_19 }; 
    wire[5:0] core_csr_decoded_decoded_lo_19 ={ core_csr_decoded_decoded_lo_hi_19 , core_csr_decoded_decoded_lo_lo_19 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_3_19 , core_csr_decoded_decoded_andMatrixInput_4_19 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_19 ={ core_csr_decoded_decoded_hi_lo_hi_19 , core_csr_decoded_decoded_andMatrixInput_5_19 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_0_19 , core_csr_decoded_decoded_andMatrixInput_1_19 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_19 ={ core_csr_decoded_decoded_hi_hi_hi_19 , core_csr_decoded_decoded_andMatrixInput_2_19 }; 
    wire[5:0] core_csr_decoded_decoded_hi_19 ={ core_csr_decoded_decoded_hi_hi_19 , core_csr_decoded_decoded_hi_lo_19 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_9_20 , core_csr_decoded_decoded_andMatrixInput_10_20 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_20 ={ core_csr_decoded_decoded_lo_lo_hi_18 , core_csr_decoded_decoded_andMatrixInput_11_18 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_6_20 , core_csr_decoded_decoded_andMatrixInput_7_20 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_20 ={ core_csr_decoded_decoded_lo_hi_hi_20 , core_csr_decoded_decoded_andMatrixInput_8_20 }; 
    wire[5:0] core_csr_decoded_decoded_lo_20 ={ core_csr_decoded_decoded_lo_hi_20 , core_csr_decoded_decoded_lo_lo_20 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_3_20 , core_csr_decoded_decoded_andMatrixInput_4_20 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_20 ={ core_csr_decoded_decoded_hi_lo_hi_20 , core_csr_decoded_decoded_andMatrixInput_5_20 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_0_20 , core_csr_decoded_decoded_andMatrixInput_1_20 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_20 ={ core_csr_decoded_decoded_hi_hi_hi_20 , core_csr_decoded_decoded_andMatrixInput_2_20 }; 
    wire[5:0] core_csr_decoded_decoded_hi_20 ={ core_csr_decoded_decoded_hi_hi_20 , core_csr_decoded_decoded_hi_lo_20 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_9_21 , core_csr_decoded_decoded_andMatrixInput_10_21 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_21 ={ core_csr_decoded_decoded_lo_lo_hi_19 , core_csr_decoded_decoded_andMatrixInput_11_19 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_6_21 , core_csr_decoded_decoded_andMatrixInput_7_21 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_21 ={ core_csr_decoded_decoded_lo_hi_hi_21 , core_csr_decoded_decoded_andMatrixInput_8_21 }; 
    wire[5:0] core_csr_decoded_decoded_lo_21 ={ core_csr_decoded_decoded_lo_hi_21 , core_csr_decoded_decoded_lo_lo_21 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_3_21 , core_csr_decoded_decoded_andMatrixInput_4_21 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_21 ={ core_csr_decoded_decoded_hi_lo_hi_21 , core_csr_decoded_decoded_andMatrixInput_5_21 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_0_21 , core_csr_decoded_decoded_andMatrixInput_1_21 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_21 ={ core_csr_decoded_decoded_hi_hi_hi_21 , core_csr_decoded_decoded_andMatrixInput_2_21 }; 
    wire[5:0] core_csr_decoded_decoded_hi_21 ={ core_csr_decoded_decoded_hi_hi_21 , core_csr_decoded_decoded_hi_lo_21 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_9_22 , core_csr_decoded_decoded_andMatrixInput_10_22 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_22 ={ core_csr_decoded_decoded_lo_lo_hi_20 , core_csr_decoded_decoded_andMatrixInput_11_20 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_6_22 , core_csr_decoded_decoded_andMatrixInput_7_22 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_22 ={ core_csr_decoded_decoded_lo_hi_hi_22 , core_csr_decoded_decoded_andMatrixInput_8_22 }; 
    wire[5:0] core_csr_decoded_decoded_lo_22 ={ core_csr_decoded_decoded_lo_hi_22 , core_csr_decoded_decoded_lo_lo_22 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_3_22 , core_csr_decoded_decoded_andMatrixInput_4_22 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_22 ={ core_csr_decoded_decoded_hi_lo_hi_22 , core_csr_decoded_decoded_andMatrixInput_5_22 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_0_22 , core_csr_decoded_decoded_andMatrixInput_1_22 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_22 ={ core_csr_decoded_decoded_hi_hi_hi_22 , core_csr_decoded_decoded_andMatrixInput_2_22 }; 
    wire[5:0] core_csr_decoded_decoded_hi_22 ={ core_csr_decoded_decoded_hi_hi_22 , core_csr_decoded_decoded_hi_lo_22 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_9_23 , core_csr_decoded_decoded_andMatrixInput_10_23 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_23 ={ core_csr_decoded_decoded_lo_lo_hi_21 , core_csr_decoded_decoded_andMatrixInput_11_21 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_6_23 , core_csr_decoded_decoded_andMatrixInput_7_23 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_23 ={ core_csr_decoded_decoded_lo_hi_hi_23 , core_csr_decoded_decoded_andMatrixInput_8_23 }; 
    wire[5:0] core_csr_decoded_decoded_lo_23 ={ core_csr_decoded_decoded_lo_hi_23 , core_csr_decoded_decoded_lo_lo_23 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_3_23 , core_csr_decoded_decoded_andMatrixInput_4_23 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_23 ={ core_csr_decoded_decoded_hi_lo_hi_23 , core_csr_decoded_decoded_andMatrixInput_5_23 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_0_23 , core_csr_decoded_decoded_andMatrixInput_1_23 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_23 ={ core_csr_decoded_decoded_hi_hi_hi_23 , core_csr_decoded_decoded_andMatrixInput_2_23 }; 
    wire[5:0] core_csr_decoded_decoded_hi_23 ={ core_csr_decoded_decoded_hi_hi_23 , core_csr_decoded_decoded_hi_lo_23 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_9_24 , core_csr_decoded_decoded_andMatrixInput_10_24 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_24 ={ core_csr_decoded_decoded_lo_lo_hi_22 , core_csr_decoded_decoded_andMatrixInput_11_22 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_6_24 , core_csr_decoded_decoded_andMatrixInput_7_24 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_24 ={ core_csr_decoded_decoded_lo_hi_hi_24 , core_csr_decoded_decoded_andMatrixInput_8_24 }; 
    wire[5:0] core_csr_decoded_decoded_lo_24 ={ core_csr_decoded_decoded_lo_hi_24 , core_csr_decoded_decoded_lo_lo_24 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_3_24 , core_csr_decoded_decoded_andMatrixInput_4_24 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_24 ={ core_csr_decoded_decoded_hi_lo_hi_24 , core_csr_decoded_decoded_andMatrixInput_5_24 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_0_24 , core_csr_decoded_decoded_andMatrixInput_1_24 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_24 ={ core_csr_decoded_decoded_hi_hi_hi_24 , core_csr_decoded_decoded_andMatrixInput_2_24 }; 
    wire[5:0] core_csr_decoded_decoded_hi_24 ={ core_csr_decoded_decoded_hi_hi_24 , core_csr_decoded_decoded_hi_lo_24 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_9_25 , core_csr_decoded_decoded_andMatrixInput_10_25 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_25 ={ core_csr_decoded_decoded_lo_lo_hi_23 , core_csr_decoded_decoded_andMatrixInput_11_23 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_6_25 , core_csr_decoded_decoded_andMatrixInput_7_25 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_25 ={ core_csr_decoded_decoded_lo_hi_hi_25 , core_csr_decoded_decoded_andMatrixInput_8_25 }; 
    wire[5:0] core_csr_decoded_decoded_lo_25 ={ core_csr_decoded_decoded_lo_hi_25 , core_csr_decoded_decoded_lo_lo_25 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_3_25 , core_csr_decoded_decoded_andMatrixInput_4_25 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_25 ={ core_csr_decoded_decoded_hi_lo_hi_25 , core_csr_decoded_decoded_andMatrixInput_5_25 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_0_25 , core_csr_decoded_decoded_andMatrixInput_1_25 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_25 ={ core_csr_decoded_decoded_hi_hi_hi_25 , core_csr_decoded_decoded_andMatrixInput_2_25 }; 
    wire[5:0] core_csr_decoded_decoded_hi_25 ={ core_csr_decoded_decoded_hi_hi_25 , core_csr_decoded_decoded_hi_lo_25 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_9_26 , core_csr_decoded_decoded_andMatrixInput_10_26 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_26 ={ core_csr_decoded_decoded_lo_lo_hi_24 , core_csr_decoded_decoded_andMatrixInput_11_24 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_6_26 , core_csr_decoded_decoded_andMatrixInput_7_26 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_26 ={ core_csr_decoded_decoded_lo_hi_hi_26 , core_csr_decoded_decoded_andMatrixInput_8_26 }; 
    wire[5:0] core_csr_decoded_decoded_lo_26 ={ core_csr_decoded_decoded_lo_hi_26 , core_csr_decoded_decoded_lo_lo_26 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_3_26 , core_csr_decoded_decoded_andMatrixInput_4_26 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_26 ={ core_csr_decoded_decoded_hi_lo_hi_26 , core_csr_decoded_decoded_andMatrixInput_5_26 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_0_26 , core_csr_decoded_decoded_andMatrixInput_1_26 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_26 ={ core_csr_decoded_decoded_hi_hi_hi_26 , core_csr_decoded_decoded_andMatrixInput_2_26 }; 
    wire[5:0] core_csr_decoded_decoded_hi_26 ={ core_csr_decoded_decoded_hi_hi_26 , core_csr_decoded_decoded_hi_lo_26 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_9_27 , core_csr_decoded_decoded_andMatrixInput_10_27 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_27 ={ core_csr_decoded_decoded_lo_lo_hi_25 , core_csr_decoded_decoded_andMatrixInput_11_25 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_6_27 , core_csr_decoded_decoded_andMatrixInput_7_27 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_27 ={ core_csr_decoded_decoded_lo_hi_hi_27 , core_csr_decoded_decoded_andMatrixInput_8_27 }; 
    wire[5:0] core_csr_decoded_decoded_lo_27 ={ core_csr_decoded_decoded_lo_hi_27 , core_csr_decoded_decoded_lo_lo_27 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_3_27 , core_csr_decoded_decoded_andMatrixInput_4_27 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_27 ={ core_csr_decoded_decoded_hi_lo_hi_27 , core_csr_decoded_decoded_andMatrixInput_5_27 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_0_27 , core_csr_decoded_decoded_andMatrixInput_1_27 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_27 ={ core_csr_decoded_decoded_hi_hi_hi_27 , core_csr_decoded_decoded_andMatrixInput_2_27 }; 
    wire[5:0] core_csr_decoded_decoded_hi_27 ={ core_csr_decoded_decoded_hi_hi_27 , core_csr_decoded_decoded_hi_lo_27 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_9_28 , core_csr_decoded_decoded_andMatrixInput_10_28 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_28 ={ core_csr_decoded_decoded_lo_lo_hi_26 , core_csr_decoded_decoded_andMatrixInput_11_26 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_6_28 , core_csr_decoded_decoded_andMatrixInput_7_28 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_28 ={ core_csr_decoded_decoded_lo_hi_hi_28 , core_csr_decoded_decoded_andMatrixInput_8_28 }; 
    wire[5:0] core_csr_decoded_decoded_lo_28 ={ core_csr_decoded_decoded_lo_hi_28 , core_csr_decoded_decoded_lo_lo_28 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_3_28 , core_csr_decoded_decoded_andMatrixInput_4_28 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_28 ={ core_csr_decoded_decoded_hi_lo_hi_28 , core_csr_decoded_decoded_andMatrixInput_5_28 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_0_28 , core_csr_decoded_decoded_andMatrixInput_1_28 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_28 ={ core_csr_decoded_decoded_hi_hi_hi_28 , core_csr_decoded_decoded_andMatrixInput_2_28 }; 
    wire[5:0] core_csr_decoded_decoded_hi_28 ={ core_csr_decoded_decoded_hi_hi_28 , core_csr_decoded_decoded_hi_lo_28 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_9_29 , core_csr_decoded_decoded_andMatrixInput_10_29 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_29 ={ core_csr_decoded_decoded_lo_lo_hi_27 , core_csr_decoded_decoded_andMatrixInput_11_27 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_6_29 , core_csr_decoded_decoded_andMatrixInput_7_29 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_29 ={ core_csr_decoded_decoded_lo_hi_hi_29 , core_csr_decoded_decoded_andMatrixInput_8_29 }; 
    wire[5:0] core_csr_decoded_decoded_lo_29 ={ core_csr_decoded_decoded_lo_hi_29 , core_csr_decoded_decoded_lo_lo_29 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_3_29 , core_csr_decoded_decoded_andMatrixInput_4_29 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_29 ={ core_csr_decoded_decoded_hi_lo_hi_29 , core_csr_decoded_decoded_andMatrixInput_5_29 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_0_29 , core_csr_decoded_decoded_andMatrixInput_1_29 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_29 ={ core_csr_decoded_decoded_hi_hi_hi_29 , core_csr_decoded_decoded_andMatrixInput_2_29 }; 
    wire[5:0] core_csr_decoded_decoded_hi_29 ={ core_csr_decoded_decoded_hi_hi_29 , core_csr_decoded_decoded_hi_lo_29 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_9_30 , core_csr_decoded_decoded_andMatrixInput_10_30 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_30 ={ core_csr_decoded_decoded_lo_lo_hi_28 , core_csr_decoded_decoded_andMatrixInput_11_28 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_6_30 , core_csr_decoded_decoded_andMatrixInput_7_30 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_30 ={ core_csr_decoded_decoded_lo_hi_hi_30 , core_csr_decoded_decoded_andMatrixInput_8_30 }; 
    wire[5:0] core_csr_decoded_decoded_lo_30 ={ core_csr_decoded_decoded_lo_hi_30 , core_csr_decoded_decoded_lo_lo_30 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_3_30 , core_csr_decoded_decoded_andMatrixInput_4_30 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_30 ={ core_csr_decoded_decoded_hi_lo_hi_30 , core_csr_decoded_decoded_andMatrixInput_5_30 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_0_30 , core_csr_decoded_decoded_andMatrixInput_1_30 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_30 ={ core_csr_decoded_decoded_hi_hi_hi_30 , core_csr_decoded_decoded_andMatrixInput_2_30 }; 
    wire[5:0] core_csr_decoded_decoded_hi_30 ={ core_csr_decoded_decoded_hi_hi_30 , core_csr_decoded_decoded_hi_lo_30 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_9_31 , core_csr_decoded_decoded_andMatrixInput_10_31 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_31 ={ core_csr_decoded_decoded_lo_lo_hi_29 , core_csr_decoded_decoded_andMatrixInput_11_29 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_6_31 , core_csr_decoded_decoded_andMatrixInput_7_31 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_31 ={ core_csr_decoded_decoded_lo_hi_hi_31 , core_csr_decoded_decoded_andMatrixInput_8_31 }; 
    wire[5:0] core_csr_decoded_decoded_lo_31 ={ core_csr_decoded_decoded_lo_hi_31 , core_csr_decoded_decoded_lo_lo_31 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_3_31 , core_csr_decoded_decoded_andMatrixInput_4_31 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_31 ={ core_csr_decoded_decoded_hi_lo_hi_31 , core_csr_decoded_decoded_andMatrixInput_5_31 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_0_31 , core_csr_decoded_decoded_andMatrixInput_1_31 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_31 ={ core_csr_decoded_decoded_hi_hi_hi_31 , core_csr_decoded_decoded_andMatrixInput_2_31 }; 
    wire[5:0] core_csr_decoded_decoded_hi_31 ={ core_csr_decoded_decoded_hi_hi_31 , core_csr_decoded_decoded_hi_lo_31 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_9_32 , core_csr_decoded_decoded_andMatrixInput_10_32 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_32 ={ core_csr_decoded_decoded_lo_lo_hi_30 , core_csr_decoded_decoded_andMatrixInput_11_30 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_6_32 , core_csr_decoded_decoded_andMatrixInput_7_32 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_32 ={ core_csr_decoded_decoded_lo_hi_hi_32 , core_csr_decoded_decoded_andMatrixInput_8_32 }; 
    wire[5:0] core_csr_decoded_decoded_lo_32 ={ core_csr_decoded_decoded_lo_hi_32 , core_csr_decoded_decoded_lo_lo_32 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_3_32 , core_csr_decoded_decoded_andMatrixInput_4_32 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_32 ={ core_csr_decoded_decoded_hi_lo_hi_32 , core_csr_decoded_decoded_andMatrixInput_5_32 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_0_32 , core_csr_decoded_decoded_andMatrixInput_1_32 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_32 ={ core_csr_decoded_decoded_hi_hi_hi_32 , core_csr_decoded_decoded_andMatrixInput_2_32 }; 
    wire[5:0] core_csr_decoded_decoded_hi_32 ={ core_csr_decoded_decoded_hi_hi_32 , core_csr_decoded_decoded_hi_lo_32 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_9_33 , core_csr_decoded_decoded_andMatrixInput_10_33 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_33 ={ core_csr_decoded_decoded_lo_lo_hi_31 , core_csr_decoded_decoded_andMatrixInput_11_31 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_6_33 , core_csr_decoded_decoded_andMatrixInput_7_33 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_33 ={ core_csr_decoded_decoded_lo_hi_hi_33 , core_csr_decoded_decoded_andMatrixInput_8_33 }; 
    wire[5:0] core_csr_decoded_decoded_lo_33 ={ core_csr_decoded_decoded_lo_hi_33 , core_csr_decoded_decoded_lo_lo_33 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_3_33 , core_csr_decoded_decoded_andMatrixInput_4_33 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_33 ={ core_csr_decoded_decoded_hi_lo_hi_33 , core_csr_decoded_decoded_andMatrixInput_5_33 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_0_33 , core_csr_decoded_decoded_andMatrixInput_1_33 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_33 ={ core_csr_decoded_decoded_hi_hi_hi_33 , core_csr_decoded_decoded_andMatrixInput_2_33 }; 
    wire[5:0] core_csr_decoded_decoded_hi_33 ={ core_csr_decoded_decoded_hi_hi_33 , core_csr_decoded_decoded_hi_lo_33 }; 
    wire core_csr_decoded_decoded_andMatrixInput_6_34 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_35 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_36 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_37 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_38 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_0_66 = core_csr_decoded_decoded_plaInput [6]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_9_34 , core_csr_decoded_decoded_andMatrixInput_10_34 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_34 ={ core_csr_decoded_decoded_lo_lo_hi_32 , core_csr_decoded_decoded_andMatrixInput_11_32 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_6_34 , core_csr_decoded_decoded_andMatrixInput_7_34 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_34 ={ core_csr_decoded_decoded_lo_hi_hi_34 , core_csr_decoded_decoded_andMatrixInput_8_34 }; 
    wire[5:0] core_csr_decoded_decoded_lo_34 ={ core_csr_decoded_decoded_lo_hi_34 , core_csr_decoded_decoded_lo_lo_34 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_3_34 , core_csr_decoded_decoded_andMatrixInput_4_34 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_34 ={ core_csr_decoded_decoded_hi_lo_hi_34 , core_csr_decoded_decoded_andMatrixInput_5_34 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_0_34 , core_csr_decoded_decoded_andMatrixInput_1_34 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_34 ={ core_csr_decoded_decoded_hi_hi_hi_34 , core_csr_decoded_decoded_andMatrixInput_2_34 }; 
    wire[5:0] core_csr_decoded_decoded_hi_34 ={ core_csr_decoded_decoded_hi_hi_34 , core_csr_decoded_decoded_hi_lo_34 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_9_35 , core_csr_decoded_decoded_andMatrixInput_10_35 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_35 ={ core_csr_decoded_decoded_lo_lo_hi_33 , core_csr_decoded_decoded_andMatrixInput_11_33 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_6_35 , core_csr_decoded_decoded_andMatrixInput_7_35 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_35 ={ core_csr_decoded_decoded_lo_hi_hi_35 , core_csr_decoded_decoded_andMatrixInput_8_35 }; 
    wire[5:0] core_csr_decoded_decoded_lo_35 ={ core_csr_decoded_decoded_lo_hi_35 , core_csr_decoded_decoded_lo_lo_35 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_3_35 , core_csr_decoded_decoded_andMatrixInput_4_35 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_35 ={ core_csr_decoded_decoded_hi_lo_hi_35 , core_csr_decoded_decoded_andMatrixInput_5_35 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_0_35 , core_csr_decoded_decoded_andMatrixInput_1_35 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_35 ={ core_csr_decoded_decoded_hi_hi_hi_35 , core_csr_decoded_decoded_andMatrixInput_2_35 }; 
    wire[5:0] core_csr_decoded_decoded_hi_35 ={ core_csr_decoded_decoded_hi_hi_35 , core_csr_decoded_decoded_hi_lo_35 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_9_36 , core_csr_decoded_decoded_andMatrixInput_10_36 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_36 ={ core_csr_decoded_decoded_lo_lo_hi_34 , core_csr_decoded_decoded_andMatrixInput_11_34 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_6_36 , core_csr_decoded_decoded_andMatrixInput_7_36 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_36 ={ core_csr_decoded_decoded_lo_hi_hi_36 , core_csr_decoded_decoded_andMatrixInput_8_36 }; 
    wire[5:0] core_csr_decoded_decoded_lo_36 ={ core_csr_decoded_decoded_lo_hi_36 , core_csr_decoded_decoded_lo_lo_36 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_3_36 , core_csr_decoded_decoded_andMatrixInput_4_36 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_36 ={ core_csr_decoded_decoded_hi_lo_hi_36 , core_csr_decoded_decoded_andMatrixInput_5_36 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_0_36 , core_csr_decoded_decoded_andMatrixInput_1_36 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_36 ={ core_csr_decoded_decoded_hi_hi_hi_36 , core_csr_decoded_decoded_andMatrixInput_2_36 }; 
    wire[5:0] core_csr_decoded_decoded_hi_36 ={ core_csr_decoded_decoded_hi_hi_36 , core_csr_decoded_decoded_hi_lo_36 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_9_37 , core_csr_decoded_decoded_andMatrixInput_10_37 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_37 ={ core_csr_decoded_decoded_lo_lo_hi_35 , core_csr_decoded_decoded_andMatrixInput_11_35 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_6_37 , core_csr_decoded_decoded_andMatrixInput_7_37 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_37 ={ core_csr_decoded_decoded_lo_hi_hi_37 , core_csr_decoded_decoded_andMatrixInput_8_37 }; 
    wire[5:0] core_csr_decoded_decoded_lo_37 ={ core_csr_decoded_decoded_lo_hi_37 , core_csr_decoded_decoded_lo_lo_37 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_3_37 , core_csr_decoded_decoded_andMatrixInput_4_37 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_37 ={ core_csr_decoded_decoded_hi_lo_hi_37 , core_csr_decoded_decoded_andMatrixInput_5_37 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_0_37 , core_csr_decoded_decoded_andMatrixInput_1_37 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_37 ={ core_csr_decoded_decoded_hi_hi_hi_37 , core_csr_decoded_decoded_andMatrixInput_2_37 }; 
    wire[5:0] core_csr_decoded_decoded_hi_37 ={ core_csr_decoded_decoded_hi_hi_37 , core_csr_decoded_decoded_hi_lo_37 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_38 ={ core_csr_decoded_decoded_andMatrixInput_8_38 , core_csr_decoded_decoded_andMatrixInput_9_38 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_5_38 , core_csr_decoded_decoded_andMatrixInput_6_38 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_38 ={ core_csr_decoded_decoded_lo_hi_hi_38 , core_csr_decoded_decoded_andMatrixInput_7_38 }; 
    wire[4:0] core_csr_decoded_decoded_lo_38 ={ core_csr_decoded_decoded_lo_hi_38 , core_csr_decoded_decoded_lo_lo_38 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_38 ={ core_csr_decoded_decoded_andMatrixInput_3_38 , core_csr_decoded_decoded_andMatrixInput_4_38 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_0_38 , core_csr_decoded_decoded_andMatrixInput_1_38 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_38 ={ core_csr_decoded_decoded_hi_hi_hi_38 , core_csr_decoded_decoded_andMatrixInput_2_38 }; 
    wire[4:0] core_csr_decoded_decoded_hi_38 ={ core_csr_decoded_decoded_hi_hi_38 , core_csr_decoded_decoded_hi_lo_38 }; 
    wire core_csr_decoded_decoded_andMatrixInput_7_39 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_40 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_41 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_42 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_43 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_44 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_45 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_46 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_47 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_48 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_49 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_50 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_51 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_52 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_53 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_54 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_55 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_56 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_57 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_58 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_59 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_60 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_61 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_62 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_63 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_64 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_65 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_66 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_97 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_98 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_99 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_100 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_101 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_102 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_103 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_104 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_105 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_106 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_107 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_108 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_109 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_110 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_111 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_112 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_113 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_114 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_115 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_116 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_117 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_118 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_119 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_120 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_121 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_122 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_123 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_124 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_125 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_126 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_127 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_159 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_160 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_161 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_162 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_163 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_164 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_165 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_166 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_167 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_168 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_169 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_170 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_171 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_172 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_173 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_174 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_175 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_176 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_177 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_178 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_179 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_180 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_181 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_182 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_183 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_184 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_185 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_186 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_187 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_188 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_189 = core_csr_decoded_decoded_plaInput [7]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_9_39 , core_csr_decoded_decoded_andMatrixInput_10_38 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_39 ={ core_csr_decoded_decoded_lo_lo_hi_36 , core_csr_decoded_decoded_andMatrixInput_11_36 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_6_39 , core_csr_decoded_decoded_andMatrixInput_7_39 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_39 ={ core_csr_decoded_decoded_lo_hi_hi_39 , core_csr_decoded_decoded_andMatrixInput_8_39 }; 
    wire[5:0] core_csr_decoded_decoded_lo_39 ={ core_csr_decoded_decoded_lo_hi_39 , core_csr_decoded_decoded_lo_lo_39 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_3_39 , core_csr_decoded_decoded_andMatrixInput_4_39 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_39 ={ core_csr_decoded_decoded_hi_lo_hi_38 , core_csr_decoded_decoded_andMatrixInput_5_39 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_0_39 , core_csr_decoded_decoded_andMatrixInput_1_39 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_39 ={ core_csr_decoded_decoded_hi_hi_hi_39 , core_csr_decoded_decoded_andMatrixInput_2_39 }; 
    wire[5:0] core_csr_decoded_decoded_hi_39 ={ core_csr_decoded_decoded_hi_hi_39 , core_csr_decoded_decoded_hi_lo_39 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_9_40 , core_csr_decoded_decoded_andMatrixInput_10_39 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_40 ={ core_csr_decoded_decoded_lo_lo_hi_37 , core_csr_decoded_decoded_andMatrixInput_11_37 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_6_40 , core_csr_decoded_decoded_andMatrixInput_7_40 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_40 ={ core_csr_decoded_decoded_lo_hi_hi_40 , core_csr_decoded_decoded_andMatrixInput_8_40 }; 
    wire[5:0] core_csr_decoded_decoded_lo_40 ={ core_csr_decoded_decoded_lo_hi_40 , core_csr_decoded_decoded_lo_lo_40 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_3_40 , core_csr_decoded_decoded_andMatrixInput_4_40 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_40 ={ core_csr_decoded_decoded_hi_lo_hi_39 , core_csr_decoded_decoded_andMatrixInput_5_40 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_0_40 , core_csr_decoded_decoded_andMatrixInput_1_40 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_40 ={ core_csr_decoded_decoded_hi_hi_hi_40 , core_csr_decoded_decoded_andMatrixInput_2_40 }; 
    wire[5:0] core_csr_decoded_decoded_hi_40 ={ core_csr_decoded_decoded_hi_hi_40 , core_csr_decoded_decoded_hi_lo_40 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_9_41 , core_csr_decoded_decoded_andMatrixInput_10_40 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_41 ={ core_csr_decoded_decoded_lo_lo_hi_38 , core_csr_decoded_decoded_andMatrixInput_11_38 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_6_41 , core_csr_decoded_decoded_andMatrixInput_7_41 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_41 ={ core_csr_decoded_decoded_lo_hi_hi_41 , core_csr_decoded_decoded_andMatrixInput_8_41 }; 
    wire[5:0] core_csr_decoded_decoded_lo_41 ={ core_csr_decoded_decoded_lo_hi_41 , core_csr_decoded_decoded_lo_lo_41 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_3_41 , core_csr_decoded_decoded_andMatrixInput_4_41 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_41 ={ core_csr_decoded_decoded_hi_lo_hi_40 , core_csr_decoded_decoded_andMatrixInput_5_41 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_0_41 , core_csr_decoded_decoded_andMatrixInput_1_41 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_41 ={ core_csr_decoded_decoded_hi_hi_hi_41 , core_csr_decoded_decoded_andMatrixInput_2_41 }; 
    wire[5:0] core_csr_decoded_decoded_hi_41 ={ core_csr_decoded_decoded_hi_hi_41 , core_csr_decoded_decoded_hi_lo_41 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_9_42 , core_csr_decoded_decoded_andMatrixInput_10_41 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_42 ={ core_csr_decoded_decoded_lo_lo_hi_39 , core_csr_decoded_decoded_andMatrixInput_11_39 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_6_42 , core_csr_decoded_decoded_andMatrixInput_7_42 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_42 ={ core_csr_decoded_decoded_lo_hi_hi_42 , core_csr_decoded_decoded_andMatrixInput_8_42 }; 
    wire[5:0] core_csr_decoded_decoded_lo_42 ={ core_csr_decoded_decoded_lo_hi_42 , core_csr_decoded_decoded_lo_lo_42 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_3_42 , core_csr_decoded_decoded_andMatrixInput_4_42 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_42 ={ core_csr_decoded_decoded_hi_lo_hi_41 , core_csr_decoded_decoded_andMatrixInput_5_42 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_0_42 , core_csr_decoded_decoded_andMatrixInput_1_42 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_42 ={ core_csr_decoded_decoded_hi_hi_hi_42 , core_csr_decoded_decoded_andMatrixInput_2_42 }; 
    wire[5:0] core_csr_decoded_decoded_hi_42 ={ core_csr_decoded_decoded_hi_hi_42 , core_csr_decoded_decoded_hi_lo_42 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_9_43 , core_csr_decoded_decoded_andMatrixInput_10_42 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_43 ={ core_csr_decoded_decoded_lo_lo_hi_40 , core_csr_decoded_decoded_andMatrixInput_11_40 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_6_43 , core_csr_decoded_decoded_andMatrixInput_7_43 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_43 ={ core_csr_decoded_decoded_lo_hi_hi_43 , core_csr_decoded_decoded_andMatrixInput_8_43 }; 
    wire[5:0] core_csr_decoded_decoded_lo_43 ={ core_csr_decoded_decoded_lo_hi_43 , core_csr_decoded_decoded_lo_lo_43 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_3_43 , core_csr_decoded_decoded_andMatrixInput_4_43 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_43 ={ core_csr_decoded_decoded_hi_lo_hi_42 , core_csr_decoded_decoded_andMatrixInput_5_43 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_0_43 , core_csr_decoded_decoded_andMatrixInput_1_43 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_43 ={ core_csr_decoded_decoded_hi_hi_hi_43 , core_csr_decoded_decoded_andMatrixInput_2_43 }; 
    wire[5:0] core_csr_decoded_decoded_hi_43 ={ core_csr_decoded_decoded_hi_hi_43 , core_csr_decoded_decoded_hi_lo_43 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_9_44 , core_csr_decoded_decoded_andMatrixInput_10_43 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_44 ={ core_csr_decoded_decoded_lo_lo_hi_41 , core_csr_decoded_decoded_andMatrixInput_11_41 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_6_44 , core_csr_decoded_decoded_andMatrixInput_7_44 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_44 ={ core_csr_decoded_decoded_lo_hi_hi_44 , core_csr_decoded_decoded_andMatrixInput_8_44 }; 
    wire[5:0] core_csr_decoded_decoded_lo_44 ={ core_csr_decoded_decoded_lo_hi_44 , core_csr_decoded_decoded_lo_lo_44 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_3_44 , core_csr_decoded_decoded_andMatrixInput_4_44 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_44 ={ core_csr_decoded_decoded_hi_lo_hi_43 , core_csr_decoded_decoded_andMatrixInput_5_44 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_0_44 , core_csr_decoded_decoded_andMatrixInput_1_44 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_44 ={ core_csr_decoded_decoded_hi_hi_hi_44 , core_csr_decoded_decoded_andMatrixInput_2_44 }; 
    wire[5:0] core_csr_decoded_decoded_hi_44 ={ core_csr_decoded_decoded_hi_hi_44 , core_csr_decoded_decoded_hi_lo_44 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_9_45 , core_csr_decoded_decoded_andMatrixInput_10_44 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_45 ={ core_csr_decoded_decoded_lo_lo_hi_42 , core_csr_decoded_decoded_andMatrixInput_11_42 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_6_45 , core_csr_decoded_decoded_andMatrixInput_7_45 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_45 ={ core_csr_decoded_decoded_lo_hi_hi_45 , core_csr_decoded_decoded_andMatrixInput_8_45 }; 
    wire[5:0] core_csr_decoded_decoded_lo_45 ={ core_csr_decoded_decoded_lo_hi_45 , core_csr_decoded_decoded_lo_lo_45 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_3_45 , core_csr_decoded_decoded_andMatrixInput_4_45 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_45 ={ core_csr_decoded_decoded_hi_lo_hi_44 , core_csr_decoded_decoded_andMatrixInput_5_45 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_0_45 , core_csr_decoded_decoded_andMatrixInput_1_45 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_45 ={ core_csr_decoded_decoded_hi_hi_hi_45 , core_csr_decoded_decoded_andMatrixInput_2_45 }; 
    wire[5:0] core_csr_decoded_decoded_hi_45 ={ core_csr_decoded_decoded_hi_hi_45 , core_csr_decoded_decoded_hi_lo_45 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_9_46 , core_csr_decoded_decoded_andMatrixInput_10_45 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_46 ={ core_csr_decoded_decoded_lo_lo_hi_43 , core_csr_decoded_decoded_andMatrixInput_11_43 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_6_46 , core_csr_decoded_decoded_andMatrixInput_7_46 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_46 ={ core_csr_decoded_decoded_lo_hi_hi_46 , core_csr_decoded_decoded_andMatrixInput_8_46 }; 
    wire[5:0] core_csr_decoded_decoded_lo_46 ={ core_csr_decoded_decoded_lo_hi_46 , core_csr_decoded_decoded_lo_lo_46 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_3_46 , core_csr_decoded_decoded_andMatrixInput_4_46 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_46 ={ core_csr_decoded_decoded_hi_lo_hi_45 , core_csr_decoded_decoded_andMatrixInput_5_46 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_0_46 , core_csr_decoded_decoded_andMatrixInput_1_46 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_46 ={ core_csr_decoded_decoded_hi_hi_hi_46 , core_csr_decoded_decoded_andMatrixInput_2_46 }; 
    wire[5:0] core_csr_decoded_decoded_hi_46 ={ core_csr_decoded_decoded_hi_hi_46 , core_csr_decoded_decoded_hi_lo_46 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_9_47 , core_csr_decoded_decoded_andMatrixInput_10_46 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_47 ={ core_csr_decoded_decoded_lo_lo_hi_44 , core_csr_decoded_decoded_andMatrixInput_11_44 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_6_47 , core_csr_decoded_decoded_andMatrixInput_7_47 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_47 ={ core_csr_decoded_decoded_lo_hi_hi_47 , core_csr_decoded_decoded_andMatrixInput_8_47 }; 
    wire[5:0] core_csr_decoded_decoded_lo_47 ={ core_csr_decoded_decoded_lo_hi_47 , core_csr_decoded_decoded_lo_lo_47 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_3_47 , core_csr_decoded_decoded_andMatrixInput_4_47 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_47 ={ core_csr_decoded_decoded_hi_lo_hi_46 , core_csr_decoded_decoded_andMatrixInput_5_47 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_0_47 , core_csr_decoded_decoded_andMatrixInput_1_47 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_47 ={ core_csr_decoded_decoded_hi_hi_hi_47 , core_csr_decoded_decoded_andMatrixInput_2_47 }; 
    wire[5:0] core_csr_decoded_decoded_hi_47 ={ core_csr_decoded_decoded_hi_hi_47 , core_csr_decoded_decoded_hi_lo_47 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_9_48 , core_csr_decoded_decoded_andMatrixInput_10_47 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_48 ={ core_csr_decoded_decoded_lo_lo_hi_45 , core_csr_decoded_decoded_andMatrixInput_11_45 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_6_48 , core_csr_decoded_decoded_andMatrixInput_7_48 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_48 ={ core_csr_decoded_decoded_lo_hi_hi_48 , core_csr_decoded_decoded_andMatrixInput_8_48 }; 
    wire[5:0] core_csr_decoded_decoded_lo_48 ={ core_csr_decoded_decoded_lo_hi_48 , core_csr_decoded_decoded_lo_lo_48 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_3_48 , core_csr_decoded_decoded_andMatrixInput_4_48 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_48 ={ core_csr_decoded_decoded_hi_lo_hi_47 , core_csr_decoded_decoded_andMatrixInput_5_48 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_0_48 , core_csr_decoded_decoded_andMatrixInput_1_48 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_48 ={ core_csr_decoded_decoded_hi_hi_hi_48 , core_csr_decoded_decoded_andMatrixInput_2_48 }; 
    wire[5:0] core_csr_decoded_decoded_hi_48 ={ core_csr_decoded_decoded_hi_hi_48 , core_csr_decoded_decoded_hi_lo_48 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_9_49 , core_csr_decoded_decoded_andMatrixInput_10_48 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_49 ={ core_csr_decoded_decoded_lo_lo_hi_46 , core_csr_decoded_decoded_andMatrixInput_11_46 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_6_49 , core_csr_decoded_decoded_andMatrixInput_7_49 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_49 ={ core_csr_decoded_decoded_lo_hi_hi_49 , core_csr_decoded_decoded_andMatrixInput_8_49 }; 
    wire[5:0] core_csr_decoded_decoded_lo_49 ={ core_csr_decoded_decoded_lo_hi_49 , core_csr_decoded_decoded_lo_lo_49 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_3_49 , core_csr_decoded_decoded_andMatrixInput_4_49 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_49 ={ core_csr_decoded_decoded_hi_lo_hi_48 , core_csr_decoded_decoded_andMatrixInput_5_49 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_0_49 , core_csr_decoded_decoded_andMatrixInput_1_49 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_49 ={ core_csr_decoded_decoded_hi_hi_hi_49 , core_csr_decoded_decoded_andMatrixInput_2_49 }; 
    wire[5:0] core_csr_decoded_decoded_hi_49 ={ core_csr_decoded_decoded_hi_hi_49 , core_csr_decoded_decoded_hi_lo_49 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_9_50 , core_csr_decoded_decoded_andMatrixInput_10_49 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_50 ={ core_csr_decoded_decoded_lo_lo_hi_47 , core_csr_decoded_decoded_andMatrixInput_11_47 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_6_50 , core_csr_decoded_decoded_andMatrixInput_7_50 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_50 ={ core_csr_decoded_decoded_lo_hi_hi_50 , core_csr_decoded_decoded_andMatrixInput_8_50 }; 
    wire[5:0] core_csr_decoded_decoded_lo_50 ={ core_csr_decoded_decoded_lo_hi_50 , core_csr_decoded_decoded_lo_lo_50 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_3_50 , core_csr_decoded_decoded_andMatrixInput_4_50 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_50 ={ core_csr_decoded_decoded_hi_lo_hi_49 , core_csr_decoded_decoded_andMatrixInput_5_50 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_0_50 , core_csr_decoded_decoded_andMatrixInput_1_50 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_50 ={ core_csr_decoded_decoded_hi_hi_hi_50 , core_csr_decoded_decoded_andMatrixInput_2_50 }; 
    wire[5:0] core_csr_decoded_decoded_hi_50 ={ core_csr_decoded_decoded_hi_hi_50 , core_csr_decoded_decoded_hi_lo_50 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_9_51 , core_csr_decoded_decoded_andMatrixInput_10_50 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_51 ={ core_csr_decoded_decoded_lo_lo_hi_48 , core_csr_decoded_decoded_andMatrixInput_11_48 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_6_51 , core_csr_decoded_decoded_andMatrixInput_7_51 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_51 ={ core_csr_decoded_decoded_lo_hi_hi_51 , core_csr_decoded_decoded_andMatrixInput_8_51 }; 
    wire[5:0] core_csr_decoded_decoded_lo_51 ={ core_csr_decoded_decoded_lo_hi_51 , core_csr_decoded_decoded_lo_lo_51 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_3_51 , core_csr_decoded_decoded_andMatrixInput_4_51 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_51 ={ core_csr_decoded_decoded_hi_lo_hi_50 , core_csr_decoded_decoded_andMatrixInput_5_51 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_0_51 , core_csr_decoded_decoded_andMatrixInput_1_51 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_51 ={ core_csr_decoded_decoded_hi_hi_hi_51 , core_csr_decoded_decoded_andMatrixInput_2_51 }; 
    wire[5:0] core_csr_decoded_decoded_hi_51 ={ core_csr_decoded_decoded_hi_hi_51 , core_csr_decoded_decoded_hi_lo_51 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_9_52 , core_csr_decoded_decoded_andMatrixInput_10_51 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_52 ={ core_csr_decoded_decoded_lo_lo_hi_49 , core_csr_decoded_decoded_andMatrixInput_11_49 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_6_52 , core_csr_decoded_decoded_andMatrixInput_7_52 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_52 ={ core_csr_decoded_decoded_lo_hi_hi_52 , core_csr_decoded_decoded_andMatrixInput_8_52 }; 
    wire[5:0] core_csr_decoded_decoded_lo_52 ={ core_csr_decoded_decoded_lo_hi_52 , core_csr_decoded_decoded_lo_lo_52 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_3_52 , core_csr_decoded_decoded_andMatrixInput_4_52 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_52 ={ core_csr_decoded_decoded_hi_lo_hi_51 , core_csr_decoded_decoded_andMatrixInput_5_52 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_0_52 , core_csr_decoded_decoded_andMatrixInput_1_52 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_52 ={ core_csr_decoded_decoded_hi_hi_hi_52 , core_csr_decoded_decoded_andMatrixInput_2_52 }; 
    wire[5:0] core_csr_decoded_decoded_hi_52 ={ core_csr_decoded_decoded_hi_hi_52 , core_csr_decoded_decoded_hi_lo_52 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_9_53 , core_csr_decoded_decoded_andMatrixInput_10_52 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_53 ={ core_csr_decoded_decoded_lo_lo_hi_50 , core_csr_decoded_decoded_andMatrixInput_11_50 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_6_53 , core_csr_decoded_decoded_andMatrixInput_7_53 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_53 ={ core_csr_decoded_decoded_lo_hi_hi_53 , core_csr_decoded_decoded_andMatrixInput_8_53 }; 
    wire[5:0] core_csr_decoded_decoded_lo_53 ={ core_csr_decoded_decoded_lo_hi_53 , core_csr_decoded_decoded_lo_lo_53 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_3_53 , core_csr_decoded_decoded_andMatrixInput_4_53 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_53 ={ core_csr_decoded_decoded_hi_lo_hi_52 , core_csr_decoded_decoded_andMatrixInput_5_53 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_0_53 , core_csr_decoded_decoded_andMatrixInput_1_53 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_53 ={ core_csr_decoded_decoded_hi_hi_hi_53 , core_csr_decoded_decoded_andMatrixInput_2_53 }; 
    wire[5:0] core_csr_decoded_decoded_hi_53 ={ core_csr_decoded_decoded_hi_hi_53 , core_csr_decoded_decoded_hi_lo_53 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_9_54 , core_csr_decoded_decoded_andMatrixInput_10_53 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_54 ={ core_csr_decoded_decoded_lo_lo_hi_51 , core_csr_decoded_decoded_andMatrixInput_11_51 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_6_54 , core_csr_decoded_decoded_andMatrixInput_7_54 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_54 ={ core_csr_decoded_decoded_lo_hi_hi_54 , core_csr_decoded_decoded_andMatrixInput_8_54 }; 
    wire[5:0] core_csr_decoded_decoded_lo_54 ={ core_csr_decoded_decoded_lo_hi_54 , core_csr_decoded_decoded_lo_lo_54 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_3_54 , core_csr_decoded_decoded_andMatrixInput_4_54 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_54 ={ core_csr_decoded_decoded_hi_lo_hi_53 , core_csr_decoded_decoded_andMatrixInput_5_54 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_0_54 , core_csr_decoded_decoded_andMatrixInput_1_54 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_54 ={ core_csr_decoded_decoded_hi_hi_hi_54 , core_csr_decoded_decoded_andMatrixInput_2_54 }; 
    wire[5:0] core_csr_decoded_decoded_hi_54 ={ core_csr_decoded_decoded_hi_hi_54 , core_csr_decoded_decoded_hi_lo_54 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_9_55 , core_csr_decoded_decoded_andMatrixInput_10_54 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_55 ={ core_csr_decoded_decoded_lo_lo_hi_52 , core_csr_decoded_decoded_andMatrixInput_11_52 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_6_55 , core_csr_decoded_decoded_andMatrixInput_7_55 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_55 ={ core_csr_decoded_decoded_lo_hi_hi_55 , core_csr_decoded_decoded_andMatrixInput_8_55 }; 
    wire[5:0] core_csr_decoded_decoded_lo_55 ={ core_csr_decoded_decoded_lo_hi_55 , core_csr_decoded_decoded_lo_lo_55 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_3_55 , core_csr_decoded_decoded_andMatrixInput_4_55 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_55 ={ core_csr_decoded_decoded_hi_lo_hi_54 , core_csr_decoded_decoded_andMatrixInput_5_55 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_0_55 , core_csr_decoded_decoded_andMatrixInput_1_55 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_55 ={ core_csr_decoded_decoded_hi_hi_hi_55 , core_csr_decoded_decoded_andMatrixInput_2_55 }; 
    wire[5:0] core_csr_decoded_decoded_hi_55 ={ core_csr_decoded_decoded_hi_hi_55 , core_csr_decoded_decoded_hi_lo_55 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_9_56 , core_csr_decoded_decoded_andMatrixInput_10_55 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_56 ={ core_csr_decoded_decoded_lo_lo_hi_53 , core_csr_decoded_decoded_andMatrixInput_11_53 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_6_56 , core_csr_decoded_decoded_andMatrixInput_7_56 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_56 ={ core_csr_decoded_decoded_lo_hi_hi_56 , core_csr_decoded_decoded_andMatrixInput_8_56 }; 
    wire[5:0] core_csr_decoded_decoded_lo_56 ={ core_csr_decoded_decoded_lo_hi_56 , core_csr_decoded_decoded_lo_lo_56 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_3_56 , core_csr_decoded_decoded_andMatrixInput_4_56 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_56 ={ core_csr_decoded_decoded_hi_lo_hi_55 , core_csr_decoded_decoded_andMatrixInput_5_56 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_0_56 , core_csr_decoded_decoded_andMatrixInput_1_56 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_56 ={ core_csr_decoded_decoded_hi_hi_hi_56 , core_csr_decoded_decoded_andMatrixInput_2_56 }; 
    wire[5:0] core_csr_decoded_decoded_hi_56 ={ core_csr_decoded_decoded_hi_hi_56 , core_csr_decoded_decoded_hi_lo_56 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_9_57 , core_csr_decoded_decoded_andMatrixInput_10_56 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_57 ={ core_csr_decoded_decoded_lo_lo_hi_54 , core_csr_decoded_decoded_andMatrixInput_11_54 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_6_57 , core_csr_decoded_decoded_andMatrixInput_7_57 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_57 ={ core_csr_decoded_decoded_lo_hi_hi_57 , core_csr_decoded_decoded_andMatrixInput_8_57 }; 
    wire[5:0] core_csr_decoded_decoded_lo_57 ={ core_csr_decoded_decoded_lo_hi_57 , core_csr_decoded_decoded_lo_lo_57 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_3_57 , core_csr_decoded_decoded_andMatrixInput_4_57 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_57 ={ core_csr_decoded_decoded_hi_lo_hi_56 , core_csr_decoded_decoded_andMatrixInput_5_57 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_0_57 , core_csr_decoded_decoded_andMatrixInput_1_57 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_57 ={ core_csr_decoded_decoded_hi_hi_hi_57 , core_csr_decoded_decoded_andMatrixInput_2_57 }; 
    wire[5:0] core_csr_decoded_decoded_hi_57 ={ core_csr_decoded_decoded_hi_hi_57 , core_csr_decoded_decoded_hi_lo_57 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_9_58 , core_csr_decoded_decoded_andMatrixInput_10_57 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_58 ={ core_csr_decoded_decoded_lo_lo_hi_55 , core_csr_decoded_decoded_andMatrixInput_11_55 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_6_58 , core_csr_decoded_decoded_andMatrixInput_7_58 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_58 ={ core_csr_decoded_decoded_lo_hi_hi_58 , core_csr_decoded_decoded_andMatrixInput_8_58 }; 
    wire[5:0] core_csr_decoded_decoded_lo_58 ={ core_csr_decoded_decoded_lo_hi_58 , core_csr_decoded_decoded_lo_lo_58 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_3_58 , core_csr_decoded_decoded_andMatrixInput_4_58 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_58 ={ core_csr_decoded_decoded_hi_lo_hi_57 , core_csr_decoded_decoded_andMatrixInput_5_58 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_0_58 , core_csr_decoded_decoded_andMatrixInput_1_58 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_58 ={ core_csr_decoded_decoded_hi_hi_hi_58 , core_csr_decoded_decoded_andMatrixInput_2_58 }; 
    wire[5:0] core_csr_decoded_decoded_hi_58 ={ core_csr_decoded_decoded_hi_hi_58 , core_csr_decoded_decoded_hi_lo_58 }; 
    wire core_csr_decoded_decoded_andMatrixInput_10_58 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_59 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_60 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_61 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_62 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_63 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_65 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_66 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_128 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_128 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_129 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_130 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_131 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_132 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_133 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_134 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_135 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_136 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_137 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_138 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_139 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_140 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_141 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_142 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_143 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_144 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_145 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_146 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_147 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_148 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_149 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_150 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_151 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_152 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_153 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_154 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_155 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_156 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_157 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_159 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_159 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_160 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_161 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_162 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_163 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_164 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_165 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_166 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_167 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_168 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_169 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_170 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_171 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_172 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_173 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_174 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_175 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_176 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_177 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_178 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_179 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_180 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_181 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_182 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_183 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_184 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_185 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_186 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_187 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_188 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_190 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_190 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_191 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_192 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_193 = core_csr_decoded_decoded_plaInput [10]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_9_59 , core_csr_decoded_decoded_andMatrixInput_10_58 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_59 ={ core_csr_decoded_decoded_lo_lo_hi_56 , core_csr_decoded_decoded_andMatrixInput_11_56 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_6_59 , core_csr_decoded_decoded_andMatrixInput_7_59 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_59 ={ core_csr_decoded_decoded_lo_hi_hi_59 , core_csr_decoded_decoded_andMatrixInput_8_59 }; 
    wire[5:0] core_csr_decoded_decoded_lo_59 ={ core_csr_decoded_decoded_lo_hi_59 , core_csr_decoded_decoded_lo_lo_59 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_3_59 , core_csr_decoded_decoded_andMatrixInput_4_59 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_59 ={ core_csr_decoded_decoded_hi_lo_hi_58 , core_csr_decoded_decoded_andMatrixInput_5_59 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_0_59 , core_csr_decoded_decoded_andMatrixInput_1_59 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_59 ={ core_csr_decoded_decoded_hi_hi_hi_59 , core_csr_decoded_decoded_andMatrixInput_2_59 }; 
    wire[5:0] core_csr_decoded_decoded_hi_59 ={ core_csr_decoded_decoded_hi_hi_59 , core_csr_decoded_decoded_hi_lo_59 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_9_60 , core_csr_decoded_decoded_andMatrixInput_10_59 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_60 ={ core_csr_decoded_decoded_lo_lo_hi_57 , core_csr_decoded_decoded_andMatrixInput_11_57 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_6_60 , core_csr_decoded_decoded_andMatrixInput_7_60 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_60 ={ core_csr_decoded_decoded_lo_hi_hi_60 , core_csr_decoded_decoded_andMatrixInput_8_60 }; 
    wire[5:0] core_csr_decoded_decoded_lo_60 ={ core_csr_decoded_decoded_lo_hi_60 , core_csr_decoded_decoded_lo_lo_60 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_3_60 , core_csr_decoded_decoded_andMatrixInput_4_60 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_60 ={ core_csr_decoded_decoded_hi_lo_hi_59 , core_csr_decoded_decoded_andMatrixInput_5_60 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_0_60 , core_csr_decoded_decoded_andMatrixInput_1_60 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_60 ={ core_csr_decoded_decoded_hi_hi_hi_60 , core_csr_decoded_decoded_andMatrixInput_2_60 }; 
    wire[5:0] core_csr_decoded_decoded_hi_60 ={ core_csr_decoded_decoded_hi_hi_60 , core_csr_decoded_decoded_hi_lo_60 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_9_61 , core_csr_decoded_decoded_andMatrixInput_10_60 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_61 ={ core_csr_decoded_decoded_lo_lo_hi_58 , core_csr_decoded_decoded_andMatrixInput_11_58 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_6_61 , core_csr_decoded_decoded_andMatrixInput_7_61 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_61 ={ core_csr_decoded_decoded_lo_hi_hi_61 , core_csr_decoded_decoded_andMatrixInput_8_61 }; 
    wire[5:0] core_csr_decoded_decoded_lo_61 ={ core_csr_decoded_decoded_lo_hi_61 , core_csr_decoded_decoded_lo_lo_61 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_3_61 , core_csr_decoded_decoded_andMatrixInput_4_61 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_61 ={ core_csr_decoded_decoded_hi_lo_hi_60 , core_csr_decoded_decoded_andMatrixInput_5_61 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_0_61 , core_csr_decoded_decoded_andMatrixInput_1_61 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_61 ={ core_csr_decoded_decoded_hi_hi_hi_61 , core_csr_decoded_decoded_andMatrixInput_2_61 }; 
    wire[5:0] core_csr_decoded_decoded_hi_61 ={ core_csr_decoded_decoded_hi_hi_61 , core_csr_decoded_decoded_hi_lo_61 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_9_62 , core_csr_decoded_decoded_andMatrixInput_10_61 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_62 ={ core_csr_decoded_decoded_lo_lo_hi_59 , core_csr_decoded_decoded_andMatrixInput_11_59 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_6_62 , core_csr_decoded_decoded_andMatrixInput_7_62 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_62 ={ core_csr_decoded_decoded_lo_hi_hi_62 , core_csr_decoded_decoded_andMatrixInput_8_62 }; 
    wire[5:0] core_csr_decoded_decoded_lo_62 ={ core_csr_decoded_decoded_lo_hi_62 , core_csr_decoded_decoded_lo_lo_62 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_3_62 , core_csr_decoded_decoded_andMatrixInput_4_62 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_62 ={ core_csr_decoded_decoded_hi_lo_hi_61 , core_csr_decoded_decoded_andMatrixInput_5_62 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_0_62 , core_csr_decoded_decoded_andMatrixInput_1_62 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_62 ={ core_csr_decoded_decoded_hi_hi_hi_62 , core_csr_decoded_decoded_andMatrixInput_2_62 }; 
    wire[5:0] core_csr_decoded_decoded_hi_62 ={ core_csr_decoded_decoded_hi_hi_62 , core_csr_decoded_decoded_hi_lo_62 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_9_63 , core_csr_decoded_decoded_andMatrixInput_10_62 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_63 ={ core_csr_decoded_decoded_lo_lo_hi_60 , core_csr_decoded_decoded_andMatrixInput_11_60 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_6_63 , core_csr_decoded_decoded_andMatrixInput_7_63 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_63 ={ core_csr_decoded_decoded_lo_hi_hi_63 , core_csr_decoded_decoded_andMatrixInput_8_63 }; 
    wire[5:0] core_csr_decoded_decoded_lo_63 ={ core_csr_decoded_decoded_lo_hi_63 , core_csr_decoded_decoded_lo_lo_63 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_3_63 , core_csr_decoded_decoded_andMatrixInput_4_63 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_63 ={ core_csr_decoded_decoded_hi_lo_hi_62 , core_csr_decoded_decoded_andMatrixInput_5_63 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_0_63 , core_csr_decoded_decoded_andMatrixInput_1_63 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_63 ={ core_csr_decoded_decoded_hi_hi_hi_63 , core_csr_decoded_decoded_andMatrixInput_2_63 }; 
    wire[5:0] core_csr_decoded_decoded_hi_63 ={ core_csr_decoded_decoded_hi_hi_63 , core_csr_decoded_decoded_hi_lo_63 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_9_64 , core_csr_decoded_decoded_andMatrixInput_10_63 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_64 ={ core_csr_decoded_decoded_lo_lo_hi_61 , core_csr_decoded_decoded_andMatrixInput_11_61 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_6_64 , core_csr_decoded_decoded_andMatrixInput_7_64 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_64 ={ core_csr_decoded_decoded_lo_hi_hi_64 , core_csr_decoded_decoded_andMatrixInput_8_64 }; 
    wire[5:0] core_csr_decoded_decoded_lo_64 ={ core_csr_decoded_decoded_lo_hi_64 , core_csr_decoded_decoded_lo_lo_64 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_3_64 , core_csr_decoded_decoded_andMatrixInput_4_64 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_64 ={ core_csr_decoded_decoded_hi_lo_hi_63 , core_csr_decoded_decoded_andMatrixInput_5_64 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_0_64 , core_csr_decoded_decoded_andMatrixInput_1_64 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_64 ={ core_csr_decoded_decoded_hi_hi_hi_64 , core_csr_decoded_decoded_andMatrixInput_2_64 }; 
    wire[5:0] core_csr_decoded_decoded_hi_64 ={ core_csr_decoded_decoded_hi_hi_64 , core_csr_decoded_decoded_hi_lo_64 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_65 ={ core_csr_decoded_decoded_andMatrixInput_9_65 , core_csr_decoded_decoded_andMatrixInput_10_64 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_6_65 , core_csr_decoded_decoded_andMatrixInput_7_65 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_65 ={ core_csr_decoded_decoded_lo_hi_hi_65 , core_csr_decoded_decoded_andMatrixInput_8_65 }; 
    wire[4:0] core_csr_decoded_decoded_lo_65 ={ core_csr_decoded_decoded_lo_hi_65 , core_csr_decoded_decoded_lo_lo_65 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_3_65 , core_csr_decoded_decoded_andMatrixInput_4_65 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_65 ={ core_csr_decoded_decoded_hi_lo_hi_64 , core_csr_decoded_decoded_andMatrixInput_5_65 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_0_65 , core_csr_decoded_decoded_andMatrixInput_1_65 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_65 ={ core_csr_decoded_decoded_hi_hi_hi_65 , core_csr_decoded_decoded_andMatrixInput_2_65 }; 
    wire[5:0] core_csr_decoded_decoded_hi_65 ={ core_csr_decoded_decoded_hi_hi_65 , core_csr_decoded_decoded_hi_lo_65 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_3_66 , core_csr_decoded_decoded_andMatrixInput_4_66 }; 
    wire[2:0] core_csr_decoded_decoded_lo_66 ={ core_csr_decoded_decoded_lo_hi_66 , core_csr_decoded_decoded_andMatrixInput_5_66 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_0_66 , core_csr_decoded_decoded_andMatrixInput_1_66 }; 
    wire[2:0] core_csr_decoded_decoded_hi_66 ={ core_csr_decoded_decoded_hi_hi_66 , core_csr_decoded_decoded_andMatrixInput_2_66 }; 
    wire core_csr_decoded_decoded_andMatrixInput_10_65 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_62 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_63 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_64 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_65 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_66 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_67 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_68 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_69 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_70 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_71 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_72 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_73 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_74 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_75 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_76 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_77 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_78 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_79 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_80 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_81 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_82 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_83 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_84 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_85 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_86 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_87 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_88 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_89 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_90 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_91 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_96 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_92 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_93 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_94 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_95 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_96 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_97 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_98 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_99 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_100 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_101 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_102 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_103 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_104 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_105 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_106 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_107 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_108 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_109 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_110 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_111 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_112 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_113 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_114 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_115 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_116 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_117 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_118 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_119 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_120 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_121 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_127 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_122 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_123 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_124 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_125 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_126 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_127 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_128 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_129 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_130 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_131 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_132 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_133 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_134 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_135 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_136 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_137 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_138 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_139 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_140 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_141 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_142 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_143 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_144 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_145 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_146 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_147 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_148 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_149 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_150 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_151 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_158 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_152 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_153 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_154 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_155 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_156 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_157 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_158 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_159 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_160 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_161 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_162 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_163 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_164 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_165 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_166 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_167 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_168 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_169 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_170 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_171 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_172 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_173 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_174 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_175 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_176 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_177 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_178 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_179 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_180 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_181 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_189 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_182 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_183 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_184 = core_csr_decoded_decoded_plaInput [11]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_185 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_66 ={ core_csr_decoded_decoded_andMatrixInput_9_66 , core_csr_decoded_decoded_andMatrixInput_10_65 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_6_66 , core_csr_decoded_decoded_andMatrixInput_7_66 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_67 ={ core_csr_decoded_decoded_lo_hi_hi_66 , core_csr_decoded_decoded_andMatrixInput_8_66 }; 
    wire[4:0] core_csr_decoded_decoded_lo_67 ={ core_csr_decoded_decoded_lo_hi_67 , core_csr_decoded_decoded_lo_lo_66 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_3_67 , core_csr_decoded_decoded_andMatrixInput_4_67 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_66 ={ core_csr_decoded_decoded_hi_lo_hi_65 , core_csr_decoded_decoded_andMatrixInput_5_67 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_0_67 , core_csr_decoded_decoded_andMatrixInput_1_67 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_67 ={ core_csr_decoded_decoded_hi_hi_hi_66 , core_csr_decoded_decoded_andMatrixInput_2_67 }; 
    wire[5:0] core_csr_decoded_decoded_hi_67 ={ core_csr_decoded_decoded_hi_hi_67 , core_csr_decoded_decoded_hi_lo_66 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_9_67 , core_csr_decoded_decoded_andMatrixInput_10_66 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_67 ={ core_csr_decoded_decoded_lo_lo_hi_62 , core_csr_decoded_decoded_andMatrixInput_11_62 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_6_67 , core_csr_decoded_decoded_andMatrixInput_7_67 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_68 ={ core_csr_decoded_decoded_lo_hi_hi_67 , core_csr_decoded_decoded_andMatrixInput_8_67 }; 
    wire[5:0] core_csr_decoded_decoded_lo_68 ={ core_csr_decoded_decoded_lo_hi_68 , core_csr_decoded_decoded_lo_lo_67 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_3_68 , core_csr_decoded_decoded_andMatrixInput_4_68 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_67 ={ core_csr_decoded_decoded_hi_lo_hi_66 , core_csr_decoded_decoded_andMatrixInput_5_68 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_0_68 , core_csr_decoded_decoded_andMatrixInput_1_68 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_68 ={ core_csr_decoded_decoded_hi_hi_hi_67 , core_csr_decoded_decoded_andMatrixInput_2_68 }; 
    wire[5:0] core_csr_decoded_decoded_hi_68 ={ core_csr_decoded_decoded_hi_hi_68 , core_csr_decoded_decoded_hi_lo_67 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_9_68 , core_csr_decoded_decoded_andMatrixInput_10_67 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_68 ={ core_csr_decoded_decoded_lo_lo_hi_63 , core_csr_decoded_decoded_andMatrixInput_11_63 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_6_68 , core_csr_decoded_decoded_andMatrixInput_7_68 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_69 ={ core_csr_decoded_decoded_lo_hi_hi_68 , core_csr_decoded_decoded_andMatrixInput_8_68 }; 
    wire[5:0] core_csr_decoded_decoded_lo_69 ={ core_csr_decoded_decoded_lo_hi_69 , core_csr_decoded_decoded_lo_lo_68 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_3_69 , core_csr_decoded_decoded_andMatrixInput_4_69 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_68 ={ core_csr_decoded_decoded_hi_lo_hi_67 , core_csr_decoded_decoded_andMatrixInput_5_69 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_0_69 , core_csr_decoded_decoded_andMatrixInput_1_69 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_69 ={ core_csr_decoded_decoded_hi_hi_hi_68 , core_csr_decoded_decoded_andMatrixInput_2_69 }; 
    wire[5:0] core_csr_decoded_decoded_hi_69 ={ core_csr_decoded_decoded_hi_hi_69 , core_csr_decoded_decoded_hi_lo_68 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_9_69 , core_csr_decoded_decoded_andMatrixInput_10_68 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_69 ={ core_csr_decoded_decoded_lo_lo_hi_64 , core_csr_decoded_decoded_andMatrixInput_11_64 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_6_69 , core_csr_decoded_decoded_andMatrixInput_7_69 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_70 ={ core_csr_decoded_decoded_lo_hi_hi_69 , core_csr_decoded_decoded_andMatrixInput_8_69 }; 
    wire[5:0] core_csr_decoded_decoded_lo_70 ={ core_csr_decoded_decoded_lo_hi_70 , core_csr_decoded_decoded_lo_lo_69 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_3_70 , core_csr_decoded_decoded_andMatrixInput_4_70 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_69 ={ core_csr_decoded_decoded_hi_lo_hi_68 , core_csr_decoded_decoded_andMatrixInput_5_70 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_0_70 , core_csr_decoded_decoded_andMatrixInput_1_70 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_70 ={ core_csr_decoded_decoded_hi_hi_hi_69 , core_csr_decoded_decoded_andMatrixInput_2_70 }; 
    wire[5:0] core_csr_decoded_decoded_hi_70 ={ core_csr_decoded_decoded_hi_hi_70 , core_csr_decoded_decoded_hi_lo_69 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_9_70 , core_csr_decoded_decoded_andMatrixInput_10_69 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_70 ={ core_csr_decoded_decoded_lo_lo_hi_65 , core_csr_decoded_decoded_andMatrixInput_11_65 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_6_70 , core_csr_decoded_decoded_andMatrixInput_7_70 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_71 ={ core_csr_decoded_decoded_lo_hi_hi_70 , core_csr_decoded_decoded_andMatrixInput_8_70 }; 
    wire[5:0] core_csr_decoded_decoded_lo_71 ={ core_csr_decoded_decoded_lo_hi_71 , core_csr_decoded_decoded_lo_lo_70 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_3_71 , core_csr_decoded_decoded_andMatrixInput_4_71 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_70 ={ core_csr_decoded_decoded_hi_lo_hi_69 , core_csr_decoded_decoded_andMatrixInput_5_71 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_0_71 , core_csr_decoded_decoded_andMatrixInput_1_71 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_71 ={ core_csr_decoded_decoded_hi_hi_hi_70 , core_csr_decoded_decoded_andMatrixInput_2_71 }; 
    wire[5:0] core_csr_decoded_decoded_hi_71 ={ core_csr_decoded_decoded_hi_hi_71 , core_csr_decoded_decoded_hi_lo_70 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_9_71 , core_csr_decoded_decoded_andMatrixInput_10_70 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_71 ={ core_csr_decoded_decoded_lo_lo_hi_66 , core_csr_decoded_decoded_andMatrixInput_11_66 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_6_71 , core_csr_decoded_decoded_andMatrixInput_7_71 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_72 ={ core_csr_decoded_decoded_lo_hi_hi_71 , core_csr_decoded_decoded_andMatrixInput_8_71 }; 
    wire[5:0] core_csr_decoded_decoded_lo_72 ={ core_csr_decoded_decoded_lo_hi_72 , core_csr_decoded_decoded_lo_lo_71 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_3_72 , core_csr_decoded_decoded_andMatrixInput_4_72 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_71 ={ core_csr_decoded_decoded_hi_lo_hi_70 , core_csr_decoded_decoded_andMatrixInput_5_72 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_0_72 , core_csr_decoded_decoded_andMatrixInput_1_72 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_72 ={ core_csr_decoded_decoded_hi_hi_hi_71 , core_csr_decoded_decoded_andMatrixInput_2_72 }; 
    wire[5:0] core_csr_decoded_decoded_hi_72 ={ core_csr_decoded_decoded_hi_hi_72 , core_csr_decoded_decoded_hi_lo_71 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_9_72 , core_csr_decoded_decoded_andMatrixInput_10_71 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_72 ={ core_csr_decoded_decoded_lo_lo_hi_67 , core_csr_decoded_decoded_andMatrixInput_11_67 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_6_72 , core_csr_decoded_decoded_andMatrixInput_7_72 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_73 ={ core_csr_decoded_decoded_lo_hi_hi_72 , core_csr_decoded_decoded_andMatrixInput_8_72 }; 
    wire[5:0] core_csr_decoded_decoded_lo_73 ={ core_csr_decoded_decoded_lo_hi_73 , core_csr_decoded_decoded_lo_lo_72 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_3_73 , core_csr_decoded_decoded_andMatrixInput_4_73 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_72 ={ core_csr_decoded_decoded_hi_lo_hi_71 , core_csr_decoded_decoded_andMatrixInput_5_73 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_0_73 , core_csr_decoded_decoded_andMatrixInput_1_73 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_73 ={ core_csr_decoded_decoded_hi_hi_hi_72 , core_csr_decoded_decoded_andMatrixInput_2_73 }; 
    wire[5:0] core_csr_decoded_decoded_hi_73 ={ core_csr_decoded_decoded_hi_hi_73 , core_csr_decoded_decoded_hi_lo_72 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_9_73 , core_csr_decoded_decoded_andMatrixInput_10_72 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_73 ={ core_csr_decoded_decoded_lo_lo_hi_68 , core_csr_decoded_decoded_andMatrixInput_11_68 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_6_73 , core_csr_decoded_decoded_andMatrixInput_7_73 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_74 ={ core_csr_decoded_decoded_lo_hi_hi_73 , core_csr_decoded_decoded_andMatrixInput_8_73 }; 
    wire[5:0] core_csr_decoded_decoded_lo_74 ={ core_csr_decoded_decoded_lo_hi_74 , core_csr_decoded_decoded_lo_lo_73 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_3_74 , core_csr_decoded_decoded_andMatrixInput_4_74 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_73 ={ core_csr_decoded_decoded_hi_lo_hi_72 , core_csr_decoded_decoded_andMatrixInput_5_74 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_0_74 , core_csr_decoded_decoded_andMatrixInput_1_74 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_74 ={ core_csr_decoded_decoded_hi_hi_hi_73 , core_csr_decoded_decoded_andMatrixInput_2_74 }; 
    wire[5:0] core_csr_decoded_decoded_hi_74 ={ core_csr_decoded_decoded_hi_hi_74 , core_csr_decoded_decoded_hi_lo_73 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_9_74 , core_csr_decoded_decoded_andMatrixInput_10_73 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_74 ={ core_csr_decoded_decoded_lo_lo_hi_69 , core_csr_decoded_decoded_andMatrixInput_11_69 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_6_74 , core_csr_decoded_decoded_andMatrixInput_7_74 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_75 ={ core_csr_decoded_decoded_lo_hi_hi_74 , core_csr_decoded_decoded_andMatrixInput_8_74 }; 
    wire[5:0] core_csr_decoded_decoded_lo_75 ={ core_csr_decoded_decoded_lo_hi_75 , core_csr_decoded_decoded_lo_lo_74 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_3_75 , core_csr_decoded_decoded_andMatrixInput_4_75 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_74 ={ core_csr_decoded_decoded_hi_lo_hi_73 , core_csr_decoded_decoded_andMatrixInput_5_75 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_0_75 , core_csr_decoded_decoded_andMatrixInput_1_75 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_75 ={ core_csr_decoded_decoded_hi_hi_hi_74 , core_csr_decoded_decoded_andMatrixInput_2_75 }; 
    wire[5:0] core_csr_decoded_decoded_hi_75 ={ core_csr_decoded_decoded_hi_hi_75 , core_csr_decoded_decoded_hi_lo_74 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_9_75 , core_csr_decoded_decoded_andMatrixInput_10_74 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_75 ={ core_csr_decoded_decoded_lo_lo_hi_70 , core_csr_decoded_decoded_andMatrixInput_11_70 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_6_75 , core_csr_decoded_decoded_andMatrixInput_7_75 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_76 ={ core_csr_decoded_decoded_lo_hi_hi_75 , core_csr_decoded_decoded_andMatrixInput_8_75 }; 
    wire[5:0] core_csr_decoded_decoded_lo_76 ={ core_csr_decoded_decoded_lo_hi_76 , core_csr_decoded_decoded_lo_lo_75 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_3_76 , core_csr_decoded_decoded_andMatrixInput_4_76 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_75 ={ core_csr_decoded_decoded_hi_lo_hi_74 , core_csr_decoded_decoded_andMatrixInput_5_76 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_0_76 , core_csr_decoded_decoded_andMatrixInput_1_76 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_76 ={ core_csr_decoded_decoded_hi_hi_hi_75 , core_csr_decoded_decoded_andMatrixInput_2_76 }; 
    wire[5:0] core_csr_decoded_decoded_hi_76 ={ core_csr_decoded_decoded_hi_hi_76 , core_csr_decoded_decoded_hi_lo_75 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_9_76 , core_csr_decoded_decoded_andMatrixInput_10_75 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_76 ={ core_csr_decoded_decoded_lo_lo_hi_71 , core_csr_decoded_decoded_andMatrixInput_11_71 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_6_76 , core_csr_decoded_decoded_andMatrixInput_7_76 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_77 ={ core_csr_decoded_decoded_lo_hi_hi_76 , core_csr_decoded_decoded_andMatrixInput_8_76 }; 
    wire[5:0] core_csr_decoded_decoded_lo_77 ={ core_csr_decoded_decoded_lo_hi_77 , core_csr_decoded_decoded_lo_lo_76 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_3_77 , core_csr_decoded_decoded_andMatrixInput_4_77 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_76 ={ core_csr_decoded_decoded_hi_lo_hi_75 , core_csr_decoded_decoded_andMatrixInput_5_77 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_0_77 , core_csr_decoded_decoded_andMatrixInput_1_77 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_77 ={ core_csr_decoded_decoded_hi_hi_hi_76 , core_csr_decoded_decoded_andMatrixInput_2_77 }; 
    wire[5:0] core_csr_decoded_decoded_hi_77 ={ core_csr_decoded_decoded_hi_hi_77 , core_csr_decoded_decoded_hi_lo_76 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_9_77 , core_csr_decoded_decoded_andMatrixInput_10_76 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_77 ={ core_csr_decoded_decoded_lo_lo_hi_72 , core_csr_decoded_decoded_andMatrixInput_11_72 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_6_77 , core_csr_decoded_decoded_andMatrixInput_7_77 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_78 ={ core_csr_decoded_decoded_lo_hi_hi_77 , core_csr_decoded_decoded_andMatrixInput_8_77 }; 
    wire[5:0] core_csr_decoded_decoded_lo_78 ={ core_csr_decoded_decoded_lo_hi_78 , core_csr_decoded_decoded_lo_lo_77 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_3_78 , core_csr_decoded_decoded_andMatrixInput_4_78 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_77 ={ core_csr_decoded_decoded_hi_lo_hi_76 , core_csr_decoded_decoded_andMatrixInput_5_78 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_0_78 , core_csr_decoded_decoded_andMatrixInput_1_78 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_78 ={ core_csr_decoded_decoded_hi_hi_hi_77 , core_csr_decoded_decoded_andMatrixInput_2_78 }; 
    wire[5:0] core_csr_decoded_decoded_hi_78 ={ core_csr_decoded_decoded_hi_hi_78 , core_csr_decoded_decoded_hi_lo_77 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_9_78 , core_csr_decoded_decoded_andMatrixInput_10_77 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_78 ={ core_csr_decoded_decoded_lo_lo_hi_73 , core_csr_decoded_decoded_andMatrixInput_11_73 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_6_78 , core_csr_decoded_decoded_andMatrixInput_7_78 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_79 ={ core_csr_decoded_decoded_lo_hi_hi_78 , core_csr_decoded_decoded_andMatrixInput_8_78 }; 
    wire[5:0] core_csr_decoded_decoded_lo_79 ={ core_csr_decoded_decoded_lo_hi_79 , core_csr_decoded_decoded_lo_lo_78 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_3_79 , core_csr_decoded_decoded_andMatrixInput_4_79 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_78 ={ core_csr_decoded_decoded_hi_lo_hi_77 , core_csr_decoded_decoded_andMatrixInput_5_79 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_0_79 , core_csr_decoded_decoded_andMatrixInput_1_79 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_79 ={ core_csr_decoded_decoded_hi_hi_hi_78 , core_csr_decoded_decoded_andMatrixInput_2_79 }; 
    wire[5:0] core_csr_decoded_decoded_hi_79 ={ core_csr_decoded_decoded_hi_hi_79 , core_csr_decoded_decoded_hi_lo_78 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_9_79 , core_csr_decoded_decoded_andMatrixInput_10_78 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_79 ={ core_csr_decoded_decoded_lo_lo_hi_74 , core_csr_decoded_decoded_andMatrixInput_11_74 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_6_79 , core_csr_decoded_decoded_andMatrixInput_7_79 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_80 ={ core_csr_decoded_decoded_lo_hi_hi_79 , core_csr_decoded_decoded_andMatrixInput_8_79 }; 
    wire[5:0] core_csr_decoded_decoded_lo_80 ={ core_csr_decoded_decoded_lo_hi_80 , core_csr_decoded_decoded_lo_lo_79 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_3_80 , core_csr_decoded_decoded_andMatrixInput_4_80 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_79 ={ core_csr_decoded_decoded_hi_lo_hi_78 , core_csr_decoded_decoded_andMatrixInput_5_80 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_0_80 , core_csr_decoded_decoded_andMatrixInput_1_80 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_80 ={ core_csr_decoded_decoded_hi_hi_hi_79 , core_csr_decoded_decoded_andMatrixInput_2_80 }; 
    wire[5:0] core_csr_decoded_decoded_hi_80 ={ core_csr_decoded_decoded_hi_hi_80 , core_csr_decoded_decoded_hi_lo_79 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_9_80 , core_csr_decoded_decoded_andMatrixInput_10_79 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_80 ={ core_csr_decoded_decoded_lo_lo_hi_75 , core_csr_decoded_decoded_andMatrixInput_11_75 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_6_80 , core_csr_decoded_decoded_andMatrixInput_7_80 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_81 ={ core_csr_decoded_decoded_lo_hi_hi_80 , core_csr_decoded_decoded_andMatrixInput_8_80 }; 
    wire[5:0] core_csr_decoded_decoded_lo_81 ={ core_csr_decoded_decoded_lo_hi_81 , core_csr_decoded_decoded_lo_lo_80 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_3_81 , core_csr_decoded_decoded_andMatrixInput_4_81 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_80 ={ core_csr_decoded_decoded_hi_lo_hi_79 , core_csr_decoded_decoded_andMatrixInput_5_81 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_0_81 , core_csr_decoded_decoded_andMatrixInput_1_81 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_81 ={ core_csr_decoded_decoded_hi_hi_hi_80 , core_csr_decoded_decoded_andMatrixInput_2_81 }; 
    wire[5:0] core_csr_decoded_decoded_hi_81 ={ core_csr_decoded_decoded_hi_hi_81 , core_csr_decoded_decoded_hi_lo_80 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_9_81 , core_csr_decoded_decoded_andMatrixInput_10_80 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_81 ={ core_csr_decoded_decoded_lo_lo_hi_76 , core_csr_decoded_decoded_andMatrixInput_11_76 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_6_81 , core_csr_decoded_decoded_andMatrixInput_7_81 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_82 ={ core_csr_decoded_decoded_lo_hi_hi_81 , core_csr_decoded_decoded_andMatrixInput_8_81 }; 
    wire[5:0] core_csr_decoded_decoded_lo_82 ={ core_csr_decoded_decoded_lo_hi_82 , core_csr_decoded_decoded_lo_lo_81 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_3_82 , core_csr_decoded_decoded_andMatrixInput_4_82 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_81 ={ core_csr_decoded_decoded_hi_lo_hi_80 , core_csr_decoded_decoded_andMatrixInput_5_82 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_0_82 , core_csr_decoded_decoded_andMatrixInput_1_82 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_82 ={ core_csr_decoded_decoded_hi_hi_hi_81 , core_csr_decoded_decoded_andMatrixInput_2_82 }; 
    wire[5:0] core_csr_decoded_decoded_hi_82 ={ core_csr_decoded_decoded_hi_hi_82 , core_csr_decoded_decoded_hi_lo_81 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_9_82 , core_csr_decoded_decoded_andMatrixInput_10_81 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_82 ={ core_csr_decoded_decoded_lo_lo_hi_77 , core_csr_decoded_decoded_andMatrixInput_11_77 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_6_82 , core_csr_decoded_decoded_andMatrixInput_7_82 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_83 ={ core_csr_decoded_decoded_lo_hi_hi_82 , core_csr_decoded_decoded_andMatrixInput_8_82 }; 
    wire[5:0] core_csr_decoded_decoded_lo_83 ={ core_csr_decoded_decoded_lo_hi_83 , core_csr_decoded_decoded_lo_lo_82 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_3_83 , core_csr_decoded_decoded_andMatrixInput_4_83 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_82 ={ core_csr_decoded_decoded_hi_lo_hi_81 , core_csr_decoded_decoded_andMatrixInput_5_83 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_0_83 , core_csr_decoded_decoded_andMatrixInput_1_83 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_83 ={ core_csr_decoded_decoded_hi_hi_hi_82 , core_csr_decoded_decoded_andMatrixInput_2_83 }; 
    wire[5:0] core_csr_decoded_decoded_hi_83 ={ core_csr_decoded_decoded_hi_hi_83 , core_csr_decoded_decoded_hi_lo_82 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_9_83 , core_csr_decoded_decoded_andMatrixInput_10_82 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_83 ={ core_csr_decoded_decoded_lo_lo_hi_78 , core_csr_decoded_decoded_andMatrixInput_11_78 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_6_83 , core_csr_decoded_decoded_andMatrixInput_7_83 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_84 ={ core_csr_decoded_decoded_lo_hi_hi_83 , core_csr_decoded_decoded_andMatrixInput_8_83 }; 
    wire[5:0] core_csr_decoded_decoded_lo_84 ={ core_csr_decoded_decoded_lo_hi_84 , core_csr_decoded_decoded_lo_lo_83 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_3_84 , core_csr_decoded_decoded_andMatrixInput_4_84 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_83 ={ core_csr_decoded_decoded_hi_lo_hi_82 , core_csr_decoded_decoded_andMatrixInput_5_84 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_0_84 , core_csr_decoded_decoded_andMatrixInput_1_84 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_84 ={ core_csr_decoded_decoded_hi_hi_hi_83 , core_csr_decoded_decoded_andMatrixInput_2_84 }; 
    wire[5:0] core_csr_decoded_decoded_hi_84 ={ core_csr_decoded_decoded_hi_hi_84 , core_csr_decoded_decoded_hi_lo_83 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_9_84 , core_csr_decoded_decoded_andMatrixInput_10_83 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_84 ={ core_csr_decoded_decoded_lo_lo_hi_79 , core_csr_decoded_decoded_andMatrixInput_11_79 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_6_84 , core_csr_decoded_decoded_andMatrixInput_7_84 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_85 ={ core_csr_decoded_decoded_lo_hi_hi_84 , core_csr_decoded_decoded_andMatrixInput_8_84 }; 
    wire[5:0] core_csr_decoded_decoded_lo_85 ={ core_csr_decoded_decoded_lo_hi_85 , core_csr_decoded_decoded_lo_lo_84 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_3_85 , core_csr_decoded_decoded_andMatrixInput_4_85 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_84 ={ core_csr_decoded_decoded_hi_lo_hi_83 , core_csr_decoded_decoded_andMatrixInput_5_85 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_0_85 , core_csr_decoded_decoded_andMatrixInput_1_85 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_85 ={ core_csr_decoded_decoded_hi_hi_hi_84 , core_csr_decoded_decoded_andMatrixInput_2_85 }; 
    wire[5:0] core_csr_decoded_decoded_hi_85 ={ core_csr_decoded_decoded_hi_hi_85 , core_csr_decoded_decoded_hi_lo_84 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_9_85 , core_csr_decoded_decoded_andMatrixInput_10_84 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_85 ={ core_csr_decoded_decoded_lo_lo_hi_80 , core_csr_decoded_decoded_andMatrixInput_11_80 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_6_85 , core_csr_decoded_decoded_andMatrixInput_7_85 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_86 ={ core_csr_decoded_decoded_lo_hi_hi_85 , core_csr_decoded_decoded_andMatrixInput_8_85 }; 
    wire[5:0] core_csr_decoded_decoded_lo_86 ={ core_csr_decoded_decoded_lo_hi_86 , core_csr_decoded_decoded_lo_lo_85 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_3_86 , core_csr_decoded_decoded_andMatrixInput_4_86 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_85 ={ core_csr_decoded_decoded_hi_lo_hi_84 , core_csr_decoded_decoded_andMatrixInput_5_86 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_0_86 , core_csr_decoded_decoded_andMatrixInput_1_86 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_86 ={ core_csr_decoded_decoded_hi_hi_hi_85 , core_csr_decoded_decoded_andMatrixInput_2_86 }; 
    wire[5:0] core_csr_decoded_decoded_hi_86 ={ core_csr_decoded_decoded_hi_hi_86 , core_csr_decoded_decoded_hi_lo_85 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_9_86 , core_csr_decoded_decoded_andMatrixInput_10_85 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_86 ={ core_csr_decoded_decoded_lo_lo_hi_81 , core_csr_decoded_decoded_andMatrixInput_11_81 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_6_86 , core_csr_decoded_decoded_andMatrixInput_7_86 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_87 ={ core_csr_decoded_decoded_lo_hi_hi_86 , core_csr_decoded_decoded_andMatrixInput_8_86 }; 
    wire[5:0] core_csr_decoded_decoded_lo_87 ={ core_csr_decoded_decoded_lo_hi_87 , core_csr_decoded_decoded_lo_lo_86 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_3_87 , core_csr_decoded_decoded_andMatrixInput_4_87 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_86 ={ core_csr_decoded_decoded_hi_lo_hi_85 , core_csr_decoded_decoded_andMatrixInput_5_87 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_0_87 , core_csr_decoded_decoded_andMatrixInput_1_87 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_87 ={ core_csr_decoded_decoded_hi_hi_hi_86 , core_csr_decoded_decoded_andMatrixInput_2_87 }; 
    wire[5:0] core_csr_decoded_decoded_hi_87 ={ core_csr_decoded_decoded_hi_hi_87 , core_csr_decoded_decoded_hi_lo_86 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_9_87 , core_csr_decoded_decoded_andMatrixInput_10_86 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_87 ={ core_csr_decoded_decoded_lo_lo_hi_82 , core_csr_decoded_decoded_andMatrixInput_11_82 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_6_87 , core_csr_decoded_decoded_andMatrixInput_7_87 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_88 ={ core_csr_decoded_decoded_lo_hi_hi_87 , core_csr_decoded_decoded_andMatrixInput_8_87 }; 
    wire[5:0] core_csr_decoded_decoded_lo_88 ={ core_csr_decoded_decoded_lo_hi_88 , core_csr_decoded_decoded_lo_lo_87 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_3_88 , core_csr_decoded_decoded_andMatrixInput_4_88 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_87 ={ core_csr_decoded_decoded_hi_lo_hi_86 , core_csr_decoded_decoded_andMatrixInput_5_88 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_0_88 , core_csr_decoded_decoded_andMatrixInput_1_88 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_88 ={ core_csr_decoded_decoded_hi_hi_hi_87 , core_csr_decoded_decoded_andMatrixInput_2_88 }; 
    wire[5:0] core_csr_decoded_decoded_hi_88 ={ core_csr_decoded_decoded_hi_hi_88 , core_csr_decoded_decoded_hi_lo_87 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_9_88 , core_csr_decoded_decoded_andMatrixInput_10_87 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_88 ={ core_csr_decoded_decoded_lo_lo_hi_83 , core_csr_decoded_decoded_andMatrixInput_11_83 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_6_88 , core_csr_decoded_decoded_andMatrixInput_7_88 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_89 ={ core_csr_decoded_decoded_lo_hi_hi_88 , core_csr_decoded_decoded_andMatrixInput_8_88 }; 
    wire[5:0] core_csr_decoded_decoded_lo_89 ={ core_csr_decoded_decoded_lo_hi_89 , core_csr_decoded_decoded_lo_lo_88 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_3_89 , core_csr_decoded_decoded_andMatrixInput_4_89 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_88 ={ core_csr_decoded_decoded_hi_lo_hi_87 , core_csr_decoded_decoded_andMatrixInput_5_89 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_0_89 , core_csr_decoded_decoded_andMatrixInput_1_89 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_89 ={ core_csr_decoded_decoded_hi_hi_hi_88 , core_csr_decoded_decoded_andMatrixInput_2_89 }; 
    wire[5:0] core_csr_decoded_decoded_hi_89 ={ core_csr_decoded_decoded_hi_hi_89 , core_csr_decoded_decoded_hi_lo_88 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_9_89 , core_csr_decoded_decoded_andMatrixInput_10_88 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_89 ={ core_csr_decoded_decoded_lo_lo_hi_84 , core_csr_decoded_decoded_andMatrixInput_11_84 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_6_89 , core_csr_decoded_decoded_andMatrixInput_7_89 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_90 ={ core_csr_decoded_decoded_lo_hi_hi_89 , core_csr_decoded_decoded_andMatrixInput_8_89 }; 
    wire[5:0] core_csr_decoded_decoded_lo_90 ={ core_csr_decoded_decoded_lo_hi_90 , core_csr_decoded_decoded_lo_lo_89 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_3_90 , core_csr_decoded_decoded_andMatrixInput_4_90 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_89 ={ core_csr_decoded_decoded_hi_lo_hi_88 , core_csr_decoded_decoded_andMatrixInput_5_90 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_0_90 , core_csr_decoded_decoded_andMatrixInput_1_90 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_90 ={ core_csr_decoded_decoded_hi_hi_hi_89 , core_csr_decoded_decoded_andMatrixInput_2_90 }; 
    wire[5:0] core_csr_decoded_decoded_hi_90 ={ core_csr_decoded_decoded_hi_hi_90 , core_csr_decoded_decoded_hi_lo_89 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_9_90 , core_csr_decoded_decoded_andMatrixInput_10_89 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_90 ={ core_csr_decoded_decoded_lo_lo_hi_85 , core_csr_decoded_decoded_andMatrixInput_11_85 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_6_90 , core_csr_decoded_decoded_andMatrixInput_7_90 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_91 ={ core_csr_decoded_decoded_lo_hi_hi_90 , core_csr_decoded_decoded_andMatrixInput_8_90 }; 
    wire[5:0] core_csr_decoded_decoded_lo_91 ={ core_csr_decoded_decoded_lo_hi_91 , core_csr_decoded_decoded_lo_lo_90 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_3_91 , core_csr_decoded_decoded_andMatrixInput_4_91 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_90 ={ core_csr_decoded_decoded_hi_lo_hi_89 , core_csr_decoded_decoded_andMatrixInput_5_91 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_0_91 , core_csr_decoded_decoded_andMatrixInput_1_91 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_91 ={ core_csr_decoded_decoded_hi_hi_hi_90 , core_csr_decoded_decoded_andMatrixInput_2_91 }; 
    wire[5:0] core_csr_decoded_decoded_hi_91 ={ core_csr_decoded_decoded_hi_hi_91 , core_csr_decoded_decoded_hi_lo_90 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_9_91 , core_csr_decoded_decoded_andMatrixInput_10_90 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_91 ={ core_csr_decoded_decoded_lo_lo_hi_86 , core_csr_decoded_decoded_andMatrixInput_11_86 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_6_91 , core_csr_decoded_decoded_andMatrixInput_7_91 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_92 ={ core_csr_decoded_decoded_lo_hi_hi_91 , core_csr_decoded_decoded_andMatrixInput_8_91 }; 
    wire[5:0] core_csr_decoded_decoded_lo_92 ={ core_csr_decoded_decoded_lo_hi_92 , core_csr_decoded_decoded_lo_lo_91 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_3_92 , core_csr_decoded_decoded_andMatrixInput_4_92 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_91 ={ core_csr_decoded_decoded_hi_lo_hi_90 , core_csr_decoded_decoded_andMatrixInput_5_92 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_0_92 , core_csr_decoded_decoded_andMatrixInput_1_92 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_92 ={ core_csr_decoded_decoded_hi_hi_hi_91 , core_csr_decoded_decoded_andMatrixInput_2_92 }; 
    wire[5:0] core_csr_decoded_decoded_hi_92 ={ core_csr_decoded_decoded_hi_hi_92 , core_csr_decoded_decoded_hi_lo_91 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_9_92 , core_csr_decoded_decoded_andMatrixInput_10_91 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_92 ={ core_csr_decoded_decoded_lo_lo_hi_87 , core_csr_decoded_decoded_andMatrixInput_11_87 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_6_92 , core_csr_decoded_decoded_andMatrixInput_7_92 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_93 ={ core_csr_decoded_decoded_lo_hi_hi_92 , core_csr_decoded_decoded_andMatrixInput_8_92 }; 
    wire[5:0] core_csr_decoded_decoded_lo_93 ={ core_csr_decoded_decoded_lo_hi_93 , core_csr_decoded_decoded_lo_lo_92 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_3_93 , core_csr_decoded_decoded_andMatrixInput_4_93 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_92 ={ core_csr_decoded_decoded_hi_lo_hi_91 , core_csr_decoded_decoded_andMatrixInput_5_93 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_0_93 , core_csr_decoded_decoded_andMatrixInput_1_93 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_93 ={ core_csr_decoded_decoded_hi_hi_hi_92 , core_csr_decoded_decoded_andMatrixInput_2_93 }; 
    wire[5:0] core_csr_decoded_decoded_hi_93 ={ core_csr_decoded_decoded_hi_hi_93 , core_csr_decoded_decoded_hi_lo_92 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_9_93 , core_csr_decoded_decoded_andMatrixInput_10_92 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_93 ={ core_csr_decoded_decoded_lo_lo_hi_88 , core_csr_decoded_decoded_andMatrixInput_11_88 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_6_93 , core_csr_decoded_decoded_andMatrixInput_7_93 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_94 ={ core_csr_decoded_decoded_lo_hi_hi_93 , core_csr_decoded_decoded_andMatrixInput_8_93 }; 
    wire[5:0] core_csr_decoded_decoded_lo_94 ={ core_csr_decoded_decoded_lo_hi_94 , core_csr_decoded_decoded_lo_lo_93 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_3_94 , core_csr_decoded_decoded_andMatrixInput_4_94 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_93 ={ core_csr_decoded_decoded_hi_lo_hi_92 , core_csr_decoded_decoded_andMatrixInput_5_94 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_0_94 , core_csr_decoded_decoded_andMatrixInput_1_94 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_94 ={ core_csr_decoded_decoded_hi_hi_hi_93 , core_csr_decoded_decoded_andMatrixInput_2_94 }; 
    wire[5:0] core_csr_decoded_decoded_hi_94 ={ core_csr_decoded_decoded_hi_hi_94 , core_csr_decoded_decoded_hi_lo_93 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_9_94 , core_csr_decoded_decoded_andMatrixInput_10_93 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_94 ={ core_csr_decoded_decoded_lo_lo_hi_89 , core_csr_decoded_decoded_andMatrixInput_11_89 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_6_94 , core_csr_decoded_decoded_andMatrixInput_7_94 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_95 ={ core_csr_decoded_decoded_lo_hi_hi_94 , core_csr_decoded_decoded_andMatrixInput_8_94 }; 
    wire[5:0] core_csr_decoded_decoded_lo_95 ={ core_csr_decoded_decoded_lo_hi_95 , core_csr_decoded_decoded_lo_lo_94 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_3_95 , core_csr_decoded_decoded_andMatrixInput_4_95 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_94 ={ core_csr_decoded_decoded_hi_lo_hi_93 , core_csr_decoded_decoded_andMatrixInput_5_95 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_0_95 , core_csr_decoded_decoded_andMatrixInput_1_95 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_95 ={ core_csr_decoded_decoded_hi_hi_hi_94 , core_csr_decoded_decoded_andMatrixInput_2_95 }; 
    wire[5:0] core_csr_decoded_decoded_hi_95 ={ core_csr_decoded_decoded_hi_hi_95 , core_csr_decoded_decoded_hi_lo_94 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_9_95 , core_csr_decoded_decoded_andMatrixInput_10_94 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_95 ={ core_csr_decoded_decoded_lo_lo_hi_90 , core_csr_decoded_decoded_andMatrixInput_11_90 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_6_95 , core_csr_decoded_decoded_andMatrixInput_7_95 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_96 ={ core_csr_decoded_decoded_lo_hi_hi_95 , core_csr_decoded_decoded_andMatrixInput_8_95 }; 
    wire[5:0] core_csr_decoded_decoded_lo_96 ={ core_csr_decoded_decoded_lo_hi_96 , core_csr_decoded_decoded_lo_lo_95 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_3_96 , core_csr_decoded_decoded_andMatrixInput_4_96 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_95 ={ core_csr_decoded_decoded_hi_lo_hi_94 , core_csr_decoded_decoded_andMatrixInput_5_96 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_0_96 , core_csr_decoded_decoded_andMatrixInput_1_96 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_96 ={ core_csr_decoded_decoded_hi_hi_hi_95 , core_csr_decoded_decoded_andMatrixInput_2_96 }; 
    wire[5:0] core_csr_decoded_decoded_hi_96 ={ core_csr_decoded_decoded_hi_hi_96 , core_csr_decoded_decoded_hi_lo_95 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_9_96 , core_csr_decoded_decoded_andMatrixInput_10_95 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_96 ={ core_csr_decoded_decoded_lo_lo_hi_91 , core_csr_decoded_decoded_andMatrixInput_11_91 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_6_96 , core_csr_decoded_decoded_andMatrixInput_7_96 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_97 ={ core_csr_decoded_decoded_lo_hi_hi_96 , core_csr_decoded_decoded_andMatrixInput_8_96 }; 
    wire[5:0] core_csr_decoded_decoded_lo_97 ={ core_csr_decoded_decoded_lo_hi_97 , core_csr_decoded_decoded_lo_lo_96 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_3_97 , core_csr_decoded_decoded_andMatrixInput_4_97 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_96 ={ core_csr_decoded_decoded_hi_lo_hi_95 , core_csr_decoded_decoded_andMatrixInput_5_97 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_0_97 , core_csr_decoded_decoded_andMatrixInput_1_97 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_97 ={ core_csr_decoded_decoded_hi_hi_hi_96 , core_csr_decoded_decoded_andMatrixInput_2_97 }; 
    wire[5:0] core_csr_decoded_decoded_hi_97 ={ core_csr_decoded_decoded_hi_hi_97 , core_csr_decoded_decoded_hi_lo_96 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_97 ={ core_csr_decoded_decoded_andMatrixInput_9_97 , core_csr_decoded_decoded_andMatrixInput_10_96 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_6_97 , core_csr_decoded_decoded_andMatrixInput_7_97 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_98 ={ core_csr_decoded_decoded_lo_hi_hi_97 , core_csr_decoded_decoded_andMatrixInput_8_97 }; 
    wire[4:0] core_csr_decoded_decoded_lo_98 ={ core_csr_decoded_decoded_lo_hi_98 , core_csr_decoded_decoded_lo_lo_97 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_3_98 , core_csr_decoded_decoded_andMatrixInput_4_98 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_97 ={ core_csr_decoded_decoded_hi_lo_hi_96 , core_csr_decoded_decoded_andMatrixInput_5_98 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_0_98 , core_csr_decoded_decoded_andMatrixInput_1_98 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_98 ={ core_csr_decoded_decoded_hi_hi_hi_97 , core_csr_decoded_decoded_andMatrixInput_2_98 }; 
    wire[5:0] core_csr_decoded_decoded_hi_98 ={ core_csr_decoded_decoded_hi_hi_98 , core_csr_decoded_decoded_hi_lo_97 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_9_98 , core_csr_decoded_decoded_andMatrixInput_10_97 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_98 ={ core_csr_decoded_decoded_lo_lo_hi_92 , core_csr_decoded_decoded_andMatrixInput_11_92 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_6_98 , core_csr_decoded_decoded_andMatrixInput_7_98 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_99 ={ core_csr_decoded_decoded_lo_hi_hi_98 , core_csr_decoded_decoded_andMatrixInput_8_98 }; 
    wire[5:0] core_csr_decoded_decoded_lo_99 ={ core_csr_decoded_decoded_lo_hi_99 , core_csr_decoded_decoded_lo_lo_98 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_3_99 , core_csr_decoded_decoded_andMatrixInput_4_99 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_98 ={ core_csr_decoded_decoded_hi_lo_hi_97 , core_csr_decoded_decoded_andMatrixInput_5_99 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_0_99 , core_csr_decoded_decoded_andMatrixInput_1_99 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_99 ={ core_csr_decoded_decoded_hi_hi_hi_98 , core_csr_decoded_decoded_andMatrixInput_2_99 }; 
    wire[5:0] core_csr_decoded_decoded_hi_99 ={ core_csr_decoded_decoded_hi_hi_99 , core_csr_decoded_decoded_hi_lo_98 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_9_99 , core_csr_decoded_decoded_andMatrixInput_10_98 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_99 ={ core_csr_decoded_decoded_lo_lo_hi_93 , core_csr_decoded_decoded_andMatrixInput_11_93 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_6_99 , core_csr_decoded_decoded_andMatrixInput_7_99 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_100 ={ core_csr_decoded_decoded_lo_hi_hi_99 , core_csr_decoded_decoded_andMatrixInput_8_99 }; 
    wire[5:0] core_csr_decoded_decoded_lo_100 ={ core_csr_decoded_decoded_lo_hi_100 , core_csr_decoded_decoded_lo_lo_99 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_3_100 , core_csr_decoded_decoded_andMatrixInput_4_100 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_99 ={ core_csr_decoded_decoded_hi_lo_hi_98 , core_csr_decoded_decoded_andMatrixInput_5_100 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_0_100 , core_csr_decoded_decoded_andMatrixInput_1_100 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_100 ={ core_csr_decoded_decoded_hi_hi_hi_99 , core_csr_decoded_decoded_andMatrixInput_2_100 }; 
    wire[5:0] core_csr_decoded_decoded_hi_100 ={ core_csr_decoded_decoded_hi_hi_100 , core_csr_decoded_decoded_hi_lo_99 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_9_100 , core_csr_decoded_decoded_andMatrixInput_10_99 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_100 ={ core_csr_decoded_decoded_lo_lo_hi_94 , core_csr_decoded_decoded_andMatrixInput_11_94 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_6_100 , core_csr_decoded_decoded_andMatrixInput_7_100 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_101 ={ core_csr_decoded_decoded_lo_hi_hi_100 , core_csr_decoded_decoded_andMatrixInput_8_100 }; 
    wire[5:0] core_csr_decoded_decoded_lo_101 ={ core_csr_decoded_decoded_lo_hi_101 , core_csr_decoded_decoded_lo_lo_100 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_3_101 , core_csr_decoded_decoded_andMatrixInput_4_101 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_100 ={ core_csr_decoded_decoded_hi_lo_hi_99 , core_csr_decoded_decoded_andMatrixInput_5_101 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_0_101 , core_csr_decoded_decoded_andMatrixInput_1_101 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_101 ={ core_csr_decoded_decoded_hi_hi_hi_100 , core_csr_decoded_decoded_andMatrixInput_2_101 }; 
    wire[5:0] core_csr_decoded_decoded_hi_101 ={ core_csr_decoded_decoded_hi_hi_101 , core_csr_decoded_decoded_hi_lo_100 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_9_101 , core_csr_decoded_decoded_andMatrixInput_10_100 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_101 ={ core_csr_decoded_decoded_lo_lo_hi_95 , core_csr_decoded_decoded_andMatrixInput_11_95 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_6_101 , core_csr_decoded_decoded_andMatrixInput_7_101 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_102 ={ core_csr_decoded_decoded_lo_hi_hi_101 , core_csr_decoded_decoded_andMatrixInput_8_101 }; 
    wire[5:0] core_csr_decoded_decoded_lo_102 ={ core_csr_decoded_decoded_lo_hi_102 , core_csr_decoded_decoded_lo_lo_101 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_3_102 , core_csr_decoded_decoded_andMatrixInput_4_102 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_101 ={ core_csr_decoded_decoded_hi_lo_hi_100 , core_csr_decoded_decoded_andMatrixInput_5_102 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_0_102 , core_csr_decoded_decoded_andMatrixInput_1_102 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_102 ={ core_csr_decoded_decoded_hi_hi_hi_101 , core_csr_decoded_decoded_andMatrixInput_2_102 }; 
    wire[5:0] core_csr_decoded_decoded_hi_102 ={ core_csr_decoded_decoded_hi_hi_102 , core_csr_decoded_decoded_hi_lo_101 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_9_102 , core_csr_decoded_decoded_andMatrixInput_10_101 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_102 ={ core_csr_decoded_decoded_lo_lo_hi_96 , core_csr_decoded_decoded_andMatrixInput_11_96 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_6_102 , core_csr_decoded_decoded_andMatrixInput_7_102 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_103 ={ core_csr_decoded_decoded_lo_hi_hi_102 , core_csr_decoded_decoded_andMatrixInput_8_102 }; 
    wire[5:0] core_csr_decoded_decoded_lo_103 ={ core_csr_decoded_decoded_lo_hi_103 , core_csr_decoded_decoded_lo_lo_102 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_3_103 , core_csr_decoded_decoded_andMatrixInput_4_103 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_102 ={ core_csr_decoded_decoded_hi_lo_hi_101 , core_csr_decoded_decoded_andMatrixInput_5_103 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_0_103 , core_csr_decoded_decoded_andMatrixInput_1_103 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_103 ={ core_csr_decoded_decoded_hi_hi_hi_102 , core_csr_decoded_decoded_andMatrixInput_2_103 }; 
    wire[5:0] core_csr_decoded_decoded_hi_103 ={ core_csr_decoded_decoded_hi_hi_103 , core_csr_decoded_decoded_hi_lo_102 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_9_103 , core_csr_decoded_decoded_andMatrixInput_10_102 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_103 ={ core_csr_decoded_decoded_lo_lo_hi_97 , core_csr_decoded_decoded_andMatrixInput_11_97 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_6_103 , core_csr_decoded_decoded_andMatrixInput_7_103 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_104 ={ core_csr_decoded_decoded_lo_hi_hi_103 , core_csr_decoded_decoded_andMatrixInput_8_103 }; 
    wire[5:0] core_csr_decoded_decoded_lo_104 ={ core_csr_decoded_decoded_lo_hi_104 , core_csr_decoded_decoded_lo_lo_103 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_3_104 , core_csr_decoded_decoded_andMatrixInput_4_104 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_103 ={ core_csr_decoded_decoded_hi_lo_hi_102 , core_csr_decoded_decoded_andMatrixInput_5_104 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_0_104 , core_csr_decoded_decoded_andMatrixInput_1_104 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_104 ={ core_csr_decoded_decoded_hi_hi_hi_103 , core_csr_decoded_decoded_andMatrixInput_2_104 }; 
    wire[5:0] core_csr_decoded_decoded_hi_104 ={ core_csr_decoded_decoded_hi_hi_104 , core_csr_decoded_decoded_hi_lo_103 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_9_104 , core_csr_decoded_decoded_andMatrixInput_10_103 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_104 ={ core_csr_decoded_decoded_lo_lo_hi_98 , core_csr_decoded_decoded_andMatrixInput_11_98 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_6_104 , core_csr_decoded_decoded_andMatrixInput_7_104 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_105 ={ core_csr_decoded_decoded_lo_hi_hi_104 , core_csr_decoded_decoded_andMatrixInput_8_104 }; 
    wire[5:0] core_csr_decoded_decoded_lo_105 ={ core_csr_decoded_decoded_lo_hi_105 , core_csr_decoded_decoded_lo_lo_104 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_3_105 , core_csr_decoded_decoded_andMatrixInput_4_105 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_104 ={ core_csr_decoded_decoded_hi_lo_hi_103 , core_csr_decoded_decoded_andMatrixInput_5_105 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_0_105 , core_csr_decoded_decoded_andMatrixInput_1_105 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_105 ={ core_csr_decoded_decoded_hi_hi_hi_104 , core_csr_decoded_decoded_andMatrixInput_2_105 }; 
    wire[5:0] core_csr_decoded_decoded_hi_105 ={ core_csr_decoded_decoded_hi_hi_105 , core_csr_decoded_decoded_hi_lo_104 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_9_105 , core_csr_decoded_decoded_andMatrixInput_10_104 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_105 ={ core_csr_decoded_decoded_lo_lo_hi_99 , core_csr_decoded_decoded_andMatrixInput_11_99 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_6_105 , core_csr_decoded_decoded_andMatrixInput_7_105 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_106 ={ core_csr_decoded_decoded_lo_hi_hi_105 , core_csr_decoded_decoded_andMatrixInput_8_105 }; 
    wire[5:0] core_csr_decoded_decoded_lo_106 ={ core_csr_decoded_decoded_lo_hi_106 , core_csr_decoded_decoded_lo_lo_105 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_3_106 , core_csr_decoded_decoded_andMatrixInput_4_106 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_105 ={ core_csr_decoded_decoded_hi_lo_hi_104 , core_csr_decoded_decoded_andMatrixInput_5_106 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_0_106 , core_csr_decoded_decoded_andMatrixInput_1_106 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_106 ={ core_csr_decoded_decoded_hi_hi_hi_105 , core_csr_decoded_decoded_andMatrixInput_2_106 }; 
    wire[5:0] core_csr_decoded_decoded_hi_106 ={ core_csr_decoded_decoded_hi_hi_106 , core_csr_decoded_decoded_hi_lo_105 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_9_106 , core_csr_decoded_decoded_andMatrixInput_10_105 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_106 ={ core_csr_decoded_decoded_lo_lo_hi_100 , core_csr_decoded_decoded_andMatrixInput_11_100 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_6_106 , core_csr_decoded_decoded_andMatrixInput_7_106 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_107 ={ core_csr_decoded_decoded_lo_hi_hi_106 , core_csr_decoded_decoded_andMatrixInput_8_106 }; 
    wire[5:0] core_csr_decoded_decoded_lo_107 ={ core_csr_decoded_decoded_lo_hi_107 , core_csr_decoded_decoded_lo_lo_106 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_3_107 , core_csr_decoded_decoded_andMatrixInput_4_107 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_106 ={ core_csr_decoded_decoded_hi_lo_hi_105 , core_csr_decoded_decoded_andMatrixInput_5_107 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_0_107 , core_csr_decoded_decoded_andMatrixInput_1_107 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_107 ={ core_csr_decoded_decoded_hi_hi_hi_106 , core_csr_decoded_decoded_andMatrixInput_2_107 }; 
    wire[5:0] core_csr_decoded_decoded_hi_107 ={ core_csr_decoded_decoded_hi_hi_107 , core_csr_decoded_decoded_hi_lo_106 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_9_107 , core_csr_decoded_decoded_andMatrixInput_10_106 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_107 ={ core_csr_decoded_decoded_lo_lo_hi_101 , core_csr_decoded_decoded_andMatrixInput_11_101 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_6_107 , core_csr_decoded_decoded_andMatrixInput_7_107 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_108 ={ core_csr_decoded_decoded_lo_hi_hi_107 , core_csr_decoded_decoded_andMatrixInput_8_107 }; 
    wire[5:0] core_csr_decoded_decoded_lo_108 ={ core_csr_decoded_decoded_lo_hi_108 , core_csr_decoded_decoded_lo_lo_107 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_3_108 , core_csr_decoded_decoded_andMatrixInput_4_108 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_107 ={ core_csr_decoded_decoded_hi_lo_hi_106 , core_csr_decoded_decoded_andMatrixInput_5_108 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_0_108 , core_csr_decoded_decoded_andMatrixInput_1_108 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_108 ={ core_csr_decoded_decoded_hi_hi_hi_107 , core_csr_decoded_decoded_andMatrixInput_2_108 }; 
    wire[5:0] core_csr_decoded_decoded_hi_108 ={ core_csr_decoded_decoded_hi_hi_108 , core_csr_decoded_decoded_hi_lo_107 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_9_108 , core_csr_decoded_decoded_andMatrixInput_10_107 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_108 ={ core_csr_decoded_decoded_lo_lo_hi_102 , core_csr_decoded_decoded_andMatrixInput_11_102 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_6_108 , core_csr_decoded_decoded_andMatrixInput_7_108 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_109 ={ core_csr_decoded_decoded_lo_hi_hi_108 , core_csr_decoded_decoded_andMatrixInput_8_108 }; 
    wire[5:0] core_csr_decoded_decoded_lo_109 ={ core_csr_decoded_decoded_lo_hi_109 , core_csr_decoded_decoded_lo_lo_108 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_3_109 , core_csr_decoded_decoded_andMatrixInput_4_109 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_108 ={ core_csr_decoded_decoded_hi_lo_hi_107 , core_csr_decoded_decoded_andMatrixInput_5_109 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_0_109 , core_csr_decoded_decoded_andMatrixInput_1_109 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_109 ={ core_csr_decoded_decoded_hi_hi_hi_108 , core_csr_decoded_decoded_andMatrixInput_2_109 }; 
    wire[5:0] core_csr_decoded_decoded_hi_109 ={ core_csr_decoded_decoded_hi_hi_109 , core_csr_decoded_decoded_hi_lo_108 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_9_109 , core_csr_decoded_decoded_andMatrixInput_10_108 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_109 ={ core_csr_decoded_decoded_lo_lo_hi_103 , core_csr_decoded_decoded_andMatrixInput_11_103 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_6_109 , core_csr_decoded_decoded_andMatrixInput_7_109 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_110 ={ core_csr_decoded_decoded_lo_hi_hi_109 , core_csr_decoded_decoded_andMatrixInput_8_109 }; 
    wire[5:0] core_csr_decoded_decoded_lo_110 ={ core_csr_decoded_decoded_lo_hi_110 , core_csr_decoded_decoded_lo_lo_109 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_3_110 , core_csr_decoded_decoded_andMatrixInput_4_110 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_109 ={ core_csr_decoded_decoded_hi_lo_hi_108 , core_csr_decoded_decoded_andMatrixInput_5_110 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_0_110 , core_csr_decoded_decoded_andMatrixInput_1_110 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_110 ={ core_csr_decoded_decoded_hi_hi_hi_109 , core_csr_decoded_decoded_andMatrixInput_2_110 }; 
    wire[5:0] core_csr_decoded_decoded_hi_110 ={ core_csr_decoded_decoded_hi_hi_110 , core_csr_decoded_decoded_hi_lo_109 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_9_110 , core_csr_decoded_decoded_andMatrixInput_10_109 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_110 ={ core_csr_decoded_decoded_lo_lo_hi_104 , core_csr_decoded_decoded_andMatrixInput_11_104 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_6_110 , core_csr_decoded_decoded_andMatrixInput_7_110 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_111 ={ core_csr_decoded_decoded_lo_hi_hi_110 , core_csr_decoded_decoded_andMatrixInput_8_110 }; 
    wire[5:0] core_csr_decoded_decoded_lo_111 ={ core_csr_decoded_decoded_lo_hi_111 , core_csr_decoded_decoded_lo_lo_110 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_3_111 , core_csr_decoded_decoded_andMatrixInput_4_111 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_110 ={ core_csr_decoded_decoded_hi_lo_hi_109 , core_csr_decoded_decoded_andMatrixInput_5_111 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_0_111 , core_csr_decoded_decoded_andMatrixInput_1_111 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_111 ={ core_csr_decoded_decoded_hi_hi_hi_110 , core_csr_decoded_decoded_andMatrixInput_2_111 }; 
    wire[5:0] core_csr_decoded_decoded_hi_111 ={ core_csr_decoded_decoded_hi_hi_111 , core_csr_decoded_decoded_hi_lo_110 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_9_111 , core_csr_decoded_decoded_andMatrixInput_10_110 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_111 ={ core_csr_decoded_decoded_lo_lo_hi_105 , core_csr_decoded_decoded_andMatrixInput_11_105 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_6_111 , core_csr_decoded_decoded_andMatrixInput_7_111 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_112 ={ core_csr_decoded_decoded_lo_hi_hi_111 , core_csr_decoded_decoded_andMatrixInput_8_111 }; 
    wire[5:0] core_csr_decoded_decoded_lo_112 ={ core_csr_decoded_decoded_lo_hi_112 , core_csr_decoded_decoded_lo_lo_111 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_3_112 , core_csr_decoded_decoded_andMatrixInput_4_112 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_111 ={ core_csr_decoded_decoded_hi_lo_hi_110 , core_csr_decoded_decoded_andMatrixInput_5_112 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_0_112 , core_csr_decoded_decoded_andMatrixInput_1_112 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_112 ={ core_csr_decoded_decoded_hi_hi_hi_111 , core_csr_decoded_decoded_andMatrixInput_2_112 }; 
    wire[5:0] core_csr_decoded_decoded_hi_112 ={ core_csr_decoded_decoded_hi_hi_112 , core_csr_decoded_decoded_hi_lo_111 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_9_112 , core_csr_decoded_decoded_andMatrixInput_10_111 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_112 ={ core_csr_decoded_decoded_lo_lo_hi_106 , core_csr_decoded_decoded_andMatrixInput_11_106 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_6_112 , core_csr_decoded_decoded_andMatrixInput_7_112 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_113 ={ core_csr_decoded_decoded_lo_hi_hi_112 , core_csr_decoded_decoded_andMatrixInput_8_112 }; 
    wire[5:0] core_csr_decoded_decoded_lo_113 ={ core_csr_decoded_decoded_lo_hi_113 , core_csr_decoded_decoded_lo_lo_112 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_3_113 , core_csr_decoded_decoded_andMatrixInput_4_113 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_112 ={ core_csr_decoded_decoded_hi_lo_hi_111 , core_csr_decoded_decoded_andMatrixInput_5_113 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_0_113 , core_csr_decoded_decoded_andMatrixInput_1_113 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_113 ={ core_csr_decoded_decoded_hi_hi_hi_112 , core_csr_decoded_decoded_andMatrixInput_2_113 }; 
    wire[5:0] core_csr_decoded_decoded_hi_113 ={ core_csr_decoded_decoded_hi_hi_113 , core_csr_decoded_decoded_hi_lo_112 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_9_113 , core_csr_decoded_decoded_andMatrixInput_10_112 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_113 ={ core_csr_decoded_decoded_lo_lo_hi_107 , core_csr_decoded_decoded_andMatrixInput_11_107 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_6_113 , core_csr_decoded_decoded_andMatrixInput_7_113 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_114 ={ core_csr_decoded_decoded_lo_hi_hi_113 , core_csr_decoded_decoded_andMatrixInput_8_113 }; 
    wire[5:0] core_csr_decoded_decoded_lo_114 ={ core_csr_decoded_decoded_lo_hi_114 , core_csr_decoded_decoded_lo_lo_113 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_3_114 , core_csr_decoded_decoded_andMatrixInput_4_114 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_113 ={ core_csr_decoded_decoded_hi_lo_hi_112 , core_csr_decoded_decoded_andMatrixInput_5_114 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_0_114 , core_csr_decoded_decoded_andMatrixInput_1_114 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_114 ={ core_csr_decoded_decoded_hi_hi_hi_113 , core_csr_decoded_decoded_andMatrixInput_2_114 }; 
    wire[5:0] core_csr_decoded_decoded_hi_114 ={ core_csr_decoded_decoded_hi_hi_114 , core_csr_decoded_decoded_hi_lo_113 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_9_114 , core_csr_decoded_decoded_andMatrixInput_10_113 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_114 ={ core_csr_decoded_decoded_lo_lo_hi_108 , core_csr_decoded_decoded_andMatrixInput_11_108 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_6_114 , core_csr_decoded_decoded_andMatrixInput_7_114 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_115 ={ core_csr_decoded_decoded_lo_hi_hi_114 , core_csr_decoded_decoded_andMatrixInput_8_114 }; 
    wire[5:0] core_csr_decoded_decoded_lo_115 ={ core_csr_decoded_decoded_lo_hi_115 , core_csr_decoded_decoded_lo_lo_114 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_3_115 , core_csr_decoded_decoded_andMatrixInput_4_115 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_114 ={ core_csr_decoded_decoded_hi_lo_hi_113 , core_csr_decoded_decoded_andMatrixInput_5_115 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_0_115 , core_csr_decoded_decoded_andMatrixInput_1_115 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_115 ={ core_csr_decoded_decoded_hi_hi_hi_114 , core_csr_decoded_decoded_andMatrixInput_2_115 }; 
    wire[5:0] core_csr_decoded_decoded_hi_115 ={ core_csr_decoded_decoded_hi_hi_115 , core_csr_decoded_decoded_hi_lo_114 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_9_115 , core_csr_decoded_decoded_andMatrixInput_10_114 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_115 ={ core_csr_decoded_decoded_lo_lo_hi_109 , core_csr_decoded_decoded_andMatrixInput_11_109 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_6_115 , core_csr_decoded_decoded_andMatrixInput_7_115 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_116 ={ core_csr_decoded_decoded_lo_hi_hi_115 , core_csr_decoded_decoded_andMatrixInput_8_115 }; 
    wire[5:0] core_csr_decoded_decoded_lo_116 ={ core_csr_decoded_decoded_lo_hi_116 , core_csr_decoded_decoded_lo_lo_115 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_3_116 , core_csr_decoded_decoded_andMatrixInput_4_116 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_115 ={ core_csr_decoded_decoded_hi_lo_hi_114 , core_csr_decoded_decoded_andMatrixInput_5_116 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_0_116 , core_csr_decoded_decoded_andMatrixInput_1_116 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_116 ={ core_csr_decoded_decoded_hi_hi_hi_115 , core_csr_decoded_decoded_andMatrixInput_2_116 }; 
    wire[5:0] core_csr_decoded_decoded_hi_116 ={ core_csr_decoded_decoded_hi_hi_116 , core_csr_decoded_decoded_hi_lo_115 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_9_116 , core_csr_decoded_decoded_andMatrixInput_10_115 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_116 ={ core_csr_decoded_decoded_lo_lo_hi_110 , core_csr_decoded_decoded_andMatrixInput_11_110 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_6_116 , core_csr_decoded_decoded_andMatrixInput_7_116 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_117 ={ core_csr_decoded_decoded_lo_hi_hi_116 , core_csr_decoded_decoded_andMatrixInput_8_116 }; 
    wire[5:0] core_csr_decoded_decoded_lo_117 ={ core_csr_decoded_decoded_lo_hi_117 , core_csr_decoded_decoded_lo_lo_116 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_3_117 , core_csr_decoded_decoded_andMatrixInput_4_117 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_116 ={ core_csr_decoded_decoded_hi_lo_hi_115 , core_csr_decoded_decoded_andMatrixInput_5_117 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_0_117 , core_csr_decoded_decoded_andMatrixInput_1_117 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_117 ={ core_csr_decoded_decoded_hi_hi_hi_116 , core_csr_decoded_decoded_andMatrixInput_2_117 }; 
    wire[5:0] core_csr_decoded_decoded_hi_117 ={ core_csr_decoded_decoded_hi_hi_117 , core_csr_decoded_decoded_hi_lo_116 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_9_117 , core_csr_decoded_decoded_andMatrixInput_10_116 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_117 ={ core_csr_decoded_decoded_lo_lo_hi_111 , core_csr_decoded_decoded_andMatrixInput_11_111 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_6_117 , core_csr_decoded_decoded_andMatrixInput_7_117 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_118 ={ core_csr_decoded_decoded_lo_hi_hi_117 , core_csr_decoded_decoded_andMatrixInput_8_117 }; 
    wire[5:0] core_csr_decoded_decoded_lo_118 ={ core_csr_decoded_decoded_lo_hi_118 , core_csr_decoded_decoded_lo_lo_117 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_3_118 , core_csr_decoded_decoded_andMatrixInput_4_118 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_117 ={ core_csr_decoded_decoded_hi_lo_hi_116 , core_csr_decoded_decoded_andMatrixInput_5_118 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_0_118 , core_csr_decoded_decoded_andMatrixInput_1_118 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_118 ={ core_csr_decoded_decoded_hi_hi_hi_117 , core_csr_decoded_decoded_andMatrixInput_2_118 }; 
    wire[5:0] core_csr_decoded_decoded_hi_118 ={ core_csr_decoded_decoded_hi_hi_118 , core_csr_decoded_decoded_hi_lo_117 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_9_118 , core_csr_decoded_decoded_andMatrixInput_10_117 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_118 ={ core_csr_decoded_decoded_lo_lo_hi_112 , core_csr_decoded_decoded_andMatrixInput_11_112 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_6_118 , core_csr_decoded_decoded_andMatrixInput_7_118 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_119 ={ core_csr_decoded_decoded_lo_hi_hi_118 , core_csr_decoded_decoded_andMatrixInput_8_118 }; 
    wire[5:0] core_csr_decoded_decoded_lo_119 ={ core_csr_decoded_decoded_lo_hi_119 , core_csr_decoded_decoded_lo_lo_118 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_3_119 , core_csr_decoded_decoded_andMatrixInput_4_119 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_118 ={ core_csr_decoded_decoded_hi_lo_hi_117 , core_csr_decoded_decoded_andMatrixInput_5_119 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_0_119 , core_csr_decoded_decoded_andMatrixInput_1_119 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_119 ={ core_csr_decoded_decoded_hi_hi_hi_118 , core_csr_decoded_decoded_andMatrixInput_2_119 }; 
    wire[5:0] core_csr_decoded_decoded_hi_119 ={ core_csr_decoded_decoded_hi_hi_119 , core_csr_decoded_decoded_hi_lo_118 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_9_119 , core_csr_decoded_decoded_andMatrixInput_10_118 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_119 ={ core_csr_decoded_decoded_lo_lo_hi_113 , core_csr_decoded_decoded_andMatrixInput_11_113 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_6_119 , core_csr_decoded_decoded_andMatrixInput_7_119 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_120 ={ core_csr_decoded_decoded_lo_hi_hi_119 , core_csr_decoded_decoded_andMatrixInput_8_119 }; 
    wire[5:0] core_csr_decoded_decoded_lo_120 ={ core_csr_decoded_decoded_lo_hi_120 , core_csr_decoded_decoded_lo_lo_119 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_3_120 , core_csr_decoded_decoded_andMatrixInput_4_120 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_119 ={ core_csr_decoded_decoded_hi_lo_hi_118 , core_csr_decoded_decoded_andMatrixInput_5_120 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_0_120 , core_csr_decoded_decoded_andMatrixInput_1_120 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_120 ={ core_csr_decoded_decoded_hi_hi_hi_119 , core_csr_decoded_decoded_andMatrixInput_2_120 }; 
    wire[5:0] core_csr_decoded_decoded_hi_120 ={ core_csr_decoded_decoded_hi_hi_120 , core_csr_decoded_decoded_hi_lo_119 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_9_120 , core_csr_decoded_decoded_andMatrixInput_10_119 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_120 ={ core_csr_decoded_decoded_lo_lo_hi_114 , core_csr_decoded_decoded_andMatrixInput_11_114 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_6_120 , core_csr_decoded_decoded_andMatrixInput_7_120 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_121 ={ core_csr_decoded_decoded_lo_hi_hi_120 , core_csr_decoded_decoded_andMatrixInput_8_120 }; 
    wire[5:0] core_csr_decoded_decoded_lo_121 ={ core_csr_decoded_decoded_lo_hi_121 , core_csr_decoded_decoded_lo_lo_120 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_3_121 , core_csr_decoded_decoded_andMatrixInput_4_121 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_120 ={ core_csr_decoded_decoded_hi_lo_hi_119 , core_csr_decoded_decoded_andMatrixInput_5_121 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_0_121 , core_csr_decoded_decoded_andMatrixInput_1_121 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_121 ={ core_csr_decoded_decoded_hi_hi_hi_120 , core_csr_decoded_decoded_andMatrixInput_2_121 }; 
    wire[5:0] core_csr_decoded_decoded_hi_121 ={ core_csr_decoded_decoded_hi_hi_121 , core_csr_decoded_decoded_hi_lo_120 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_9_121 , core_csr_decoded_decoded_andMatrixInput_10_120 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_121 ={ core_csr_decoded_decoded_lo_lo_hi_115 , core_csr_decoded_decoded_andMatrixInput_11_115 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_6_121 , core_csr_decoded_decoded_andMatrixInput_7_121 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_122 ={ core_csr_decoded_decoded_lo_hi_hi_121 , core_csr_decoded_decoded_andMatrixInput_8_121 }; 
    wire[5:0] core_csr_decoded_decoded_lo_122 ={ core_csr_decoded_decoded_lo_hi_122 , core_csr_decoded_decoded_lo_lo_121 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_3_122 , core_csr_decoded_decoded_andMatrixInput_4_122 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_121 ={ core_csr_decoded_decoded_hi_lo_hi_120 , core_csr_decoded_decoded_andMatrixInput_5_122 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_0_122 , core_csr_decoded_decoded_andMatrixInput_1_122 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_122 ={ core_csr_decoded_decoded_hi_hi_hi_121 , core_csr_decoded_decoded_andMatrixInput_2_122 }; 
    wire[5:0] core_csr_decoded_decoded_hi_122 ={ core_csr_decoded_decoded_hi_hi_122 , core_csr_decoded_decoded_hi_lo_121 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_9_122 , core_csr_decoded_decoded_andMatrixInput_10_121 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_122 ={ core_csr_decoded_decoded_lo_lo_hi_116 , core_csr_decoded_decoded_andMatrixInput_11_116 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_6_122 , core_csr_decoded_decoded_andMatrixInput_7_122 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_123 ={ core_csr_decoded_decoded_lo_hi_hi_122 , core_csr_decoded_decoded_andMatrixInput_8_122 }; 
    wire[5:0] core_csr_decoded_decoded_lo_123 ={ core_csr_decoded_decoded_lo_hi_123 , core_csr_decoded_decoded_lo_lo_122 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_3_123 , core_csr_decoded_decoded_andMatrixInput_4_123 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_122 ={ core_csr_decoded_decoded_hi_lo_hi_121 , core_csr_decoded_decoded_andMatrixInput_5_123 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_0_123 , core_csr_decoded_decoded_andMatrixInput_1_123 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_123 ={ core_csr_decoded_decoded_hi_hi_hi_122 , core_csr_decoded_decoded_andMatrixInput_2_123 }; 
    wire[5:0] core_csr_decoded_decoded_hi_123 ={ core_csr_decoded_decoded_hi_hi_123 , core_csr_decoded_decoded_hi_lo_122 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_9_123 , core_csr_decoded_decoded_andMatrixInput_10_122 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_123 ={ core_csr_decoded_decoded_lo_lo_hi_117 , core_csr_decoded_decoded_andMatrixInput_11_117 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_6_123 , core_csr_decoded_decoded_andMatrixInput_7_123 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_124 ={ core_csr_decoded_decoded_lo_hi_hi_123 , core_csr_decoded_decoded_andMatrixInput_8_123 }; 
    wire[5:0] core_csr_decoded_decoded_lo_124 ={ core_csr_decoded_decoded_lo_hi_124 , core_csr_decoded_decoded_lo_lo_123 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_3_124 , core_csr_decoded_decoded_andMatrixInput_4_124 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_123 ={ core_csr_decoded_decoded_hi_lo_hi_122 , core_csr_decoded_decoded_andMatrixInput_5_124 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_0_124 , core_csr_decoded_decoded_andMatrixInput_1_124 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_124 ={ core_csr_decoded_decoded_hi_hi_hi_123 , core_csr_decoded_decoded_andMatrixInput_2_124 }; 
    wire[5:0] core_csr_decoded_decoded_hi_124 ={ core_csr_decoded_decoded_hi_hi_124 , core_csr_decoded_decoded_hi_lo_123 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_9_124 , core_csr_decoded_decoded_andMatrixInput_10_123 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_124 ={ core_csr_decoded_decoded_lo_lo_hi_118 , core_csr_decoded_decoded_andMatrixInput_11_118 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_6_124 , core_csr_decoded_decoded_andMatrixInput_7_124 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_125 ={ core_csr_decoded_decoded_lo_hi_hi_124 , core_csr_decoded_decoded_andMatrixInput_8_124 }; 
    wire[5:0] core_csr_decoded_decoded_lo_125 ={ core_csr_decoded_decoded_lo_hi_125 , core_csr_decoded_decoded_lo_lo_124 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_3_125 , core_csr_decoded_decoded_andMatrixInput_4_125 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_124 ={ core_csr_decoded_decoded_hi_lo_hi_123 , core_csr_decoded_decoded_andMatrixInput_5_125 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_0_125 , core_csr_decoded_decoded_andMatrixInput_1_125 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_125 ={ core_csr_decoded_decoded_hi_hi_hi_124 , core_csr_decoded_decoded_andMatrixInput_2_125 }; 
    wire[5:0] core_csr_decoded_decoded_hi_125 ={ core_csr_decoded_decoded_hi_hi_125 , core_csr_decoded_decoded_hi_lo_124 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_9_125 , core_csr_decoded_decoded_andMatrixInput_10_124 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_125 ={ core_csr_decoded_decoded_lo_lo_hi_119 , core_csr_decoded_decoded_andMatrixInput_11_119 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_6_125 , core_csr_decoded_decoded_andMatrixInput_7_125 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_126 ={ core_csr_decoded_decoded_lo_hi_hi_125 , core_csr_decoded_decoded_andMatrixInput_8_125 }; 
    wire[5:0] core_csr_decoded_decoded_lo_126 ={ core_csr_decoded_decoded_lo_hi_126 , core_csr_decoded_decoded_lo_lo_125 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_3_126 , core_csr_decoded_decoded_andMatrixInput_4_126 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_125 ={ core_csr_decoded_decoded_hi_lo_hi_124 , core_csr_decoded_decoded_andMatrixInput_5_126 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_0_126 , core_csr_decoded_decoded_andMatrixInput_1_126 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_126 ={ core_csr_decoded_decoded_hi_hi_hi_125 , core_csr_decoded_decoded_andMatrixInput_2_126 }; 
    wire[5:0] core_csr_decoded_decoded_hi_126 ={ core_csr_decoded_decoded_hi_hi_126 , core_csr_decoded_decoded_hi_lo_125 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_9_126 , core_csr_decoded_decoded_andMatrixInput_10_125 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_126 ={ core_csr_decoded_decoded_lo_lo_hi_120 , core_csr_decoded_decoded_andMatrixInput_11_120 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_6_126 , core_csr_decoded_decoded_andMatrixInput_7_126 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_127 ={ core_csr_decoded_decoded_lo_hi_hi_126 , core_csr_decoded_decoded_andMatrixInput_8_126 }; 
    wire[5:0] core_csr_decoded_decoded_lo_127 ={ core_csr_decoded_decoded_lo_hi_127 , core_csr_decoded_decoded_lo_lo_126 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_3_127 , core_csr_decoded_decoded_andMatrixInput_4_127 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_126 ={ core_csr_decoded_decoded_hi_lo_hi_125 , core_csr_decoded_decoded_andMatrixInput_5_127 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_0_127 , core_csr_decoded_decoded_andMatrixInput_1_127 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_127 ={ core_csr_decoded_decoded_hi_hi_hi_126 , core_csr_decoded_decoded_andMatrixInput_2_127 }; 
    wire[5:0] core_csr_decoded_decoded_hi_127 ={ core_csr_decoded_decoded_hi_hi_127 , core_csr_decoded_decoded_hi_lo_126 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_9_127 , core_csr_decoded_decoded_andMatrixInput_10_126 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_127 ={ core_csr_decoded_decoded_lo_lo_hi_121 , core_csr_decoded_decoded_andMatrixInput_11_121 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_6_127 , core_csr_decoded_decoded_andMatrixInput_7_127 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_128 ={ core_csr_decoded_decoded_lo_hi_hi_127 , core_csr_decoded_decoded_andMatrixInput_8_127 }; 
    wire[5:0] core_csr_decoded_decoded_lo_128 ={ core_csr_decoded_decoded_lo_hi_128 , core_csr_decoded_decoded_lo_lo_127 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_3_128 , core_csr_decoded_decoded_andMatrixInput_4_128 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_127 ={ core_csr_decoded_decoded_hi_lo_hi_126 , core_csr_decoded_decoded_andMatrixInput_5_128 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_0_128 , core_csr_decoded_decoded_andMatrixInput_1_128 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_128 ={ core_csr_decoded_decoded_hi_hi_hi_127 , core_csr_decoded_decoded_andMatrixInput_2_128 }; 
    wire[5:0] core_csr_decoded_decoded_hi_128 ={ core_csr_decoded_decoded_hi_hi_128 , core_csr_decoded_decoded_hi_lo_127 }; 
    wire core_csr_decoded_decoded_andMatrixInput_7_128 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_129 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_130 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_131 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_132 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_133 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_134 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_135 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_136 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_137 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_138 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_139 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_140 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_141 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_142 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_143 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_144 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_145 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_146 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_147 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_148 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_149 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_150 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_151 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_152 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_153 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_154 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_155 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_156 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_157 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_158 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_159 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_160 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_161 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_162 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_163 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_164 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_165 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_166 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_167 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_168 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_169 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_170 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_171 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_172 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_173 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_174 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_175 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_176 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_177 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_178 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_179 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_180 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_181 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_182 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_183 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_184 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_185 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_186 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_187 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_188 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_189 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_128 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_129 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_130 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_131 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_132 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_133 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_134 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_135 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_136 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_137 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_138 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_139 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_140 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_141 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_142 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_143 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_144 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_145 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_146 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_147 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_148 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_149 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_150 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_151 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_152 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_153 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_154 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_155 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_156 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_157 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_158 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_159 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_160 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_161 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_162 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_163 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_164 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_165 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_166 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_167 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_168 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_169 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_170 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_171 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_172 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_173 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_174 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_175 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_176 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_177 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_178 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_179 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_180 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_181 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_182 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_183 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_184 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_185 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_186 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_187 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_188 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_189 = core_csr_decoded_decoded_invInputs [9]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_128 ={ core_csr_decoded_decoded_andMatrixInput_9_128 , core_csr_decoded_decoded_andMatrixInput_10_127 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_6_128 , core_csr_decoded_decoded_andMatrixInput_7_128 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_129 ={ core_csr_decoded_decoded_lo_hi_hi_128 , core_csr_decoded_decoded_andMatrixInput_8_128 }; 
    wire[4:0] core_csr_decoded_decoded_lo_129 ={ core_csr_decoded_decoded_lo_hi_129 , core_csr_decoded_decoded_lo_lo_128 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_3_129 , core_csr_decoded_decoded_andMatrixInput_4_129 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_128 ={ core_csr_decoded_decoded_hi_lo_hi_127 , core_csr_decoded_decoded_andMatrixInput_5_129 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_0_129 , core_csr_decoded_decoded_andMatrixInput_1_129 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_129 ={ core_csr_decoded_decoded_hi_hi_hi_128 , core_csr_decoded_decoded_andMatrixInput_2_129 }; 
    wire[5:0] core_csr_decoded_decoded_hi_129 ={ core_csr_decoded_decoded_hi_hi_129 , core_csr_decoded_decoded_hi_lo_128 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_9_129 , core_csr_decoded_decoded_andMatrixInput_10_128 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_129 ={ core_csr_decoded_decoded_lo_lo_hi_122 , core_csr_decoded_decoded_andMatrixInput_11_122 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_6_129 , core_csr_decoded_decoded_andMatrixInput_7_129 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_130 ={ core_csr_decoded_decoded_lo_hi_hi_129 , core_csr_decoded_decoded_andMatrixInput_8_129 }; 
    wire[5:0] core_csr_decoded_decoded_lo_130 ={ core_csr_decoded_decoded_lo_hi_130 , core_csr_decoded_decoded_lo_lo_129 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_3_130 , core_csr_decoded_decoded_andMatrixInput_4_130 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_129 ={ core_csr_decoded_decoded_hi_lo_hi_128 , core_csr_decoded_decoded_andMatrixInput_5_130 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_0_130 , core_csr_decoded_decoded_andMatrixInput_1_130 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_130 ={ core_csr_decoded_decoded_hi_hi_hi_129 , core_csr_decoded_decoded_andMatrixInput_2_130 }; 
    wire[5:0] core_csr_decoded_decoded_hi_130 ={ core_csr_decoded_decoded_hi_hi_130 , core_csr_decoded_decoded_hi_lo_129 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_9_130 , core_csr_decoded_decoded_andMatrixInput_10_129 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_130 ={ core_csr_decoded_decoded_lo_lo_hi_123 , core_csr_decoded_decoded_andMatrixInput_11_123 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_130 ={ core_csr_decoded_decoded_andMatrixInput_6_130 , core_csr_decoded_decoded_andMatrixInput_7_130 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_131 ={ core_csr_decoded_decoded_lo_hi_hi_130 , core_csr_decoded_decoded_andMatrixInput_8_130 }; 
    wire[5:0] core_csr_decoded_decoded_lo_131 ={ core_csr_decoded_decoded_lo_hi_131 , core_csr_decoded_decoded_lo_lo_130 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_3_131 , core_csr_decoded_decoded_andMatrixInput_4_131 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_130 ={ core_csr_decoded_decoded_hi_lo_hi_129 , core_csr_decoded_decoded_andMatrixInput_5_131 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_130 ={ core_csr_decoded_decoded_andMatrixInput_0_131 , core_csr_decoded_decoded_andMatrixInput_1_131 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_131 ={ core_csr_decoded_decoded_hi_hi_hi_130 , core_csr_decoded_decoded_andMatrixInput_2_131 }; 
    wire[5:0] core_csr_decoded_decoded_hi_131 ={ core_csr_decoded_decoded_hi_hi_131 , core_csr_decoded_decoded_hi_lo_130 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_9_131 , core_csr_decoded_decoded_andMatrixInput_10_130 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_131 ={ core_csr_decoded_decoded_lo_lo_hi_124 , core_csr_decoded_decoded_andMatrixInput_11_124 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_131 ={ core_csr_decoded_decoded_andMatrixInput_6_131 , core_csr_decoded_decoded_andMatrixInput_7_131 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_132 ={ core_csr_decoded_decoded_lo_hi_hi_131 , core_csr_decoded_decoded_andMatrixInput_8_131 }; 
    wire[5:0] core_csr_decoded_decoded_lo_132 ={ core_csr_decoded_decoded_lo_hi_132 , core_csr_decoded_decoded_lo_lo_131 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_130 ={ core_csr_decoded_decoded_andMatrixInput_3_132 , core_csr_decoded_decoded_andMatrixInput_4_132 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_131 ={ core_csr_decoded_decoded_hi_lo_hi_130 , core_csr_decoded_decoded_andMatrixInput_5_132 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_131 ={ core_csr_decoded_decoded_andMatrixInput_0_132 , core_csr_decoded_decoded_andMatrixInput_1_132 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_132 ={ core_csr_decoded_decoded_hi_hi_hi_131 , core_csr_decoded_decoded_andMatrixInput_2_132 }; 
    wire[5:0] core_csr_decoded_decoded_hi_132 ={ core_csr_decoded_decoded_hi_hi_132 , core_csr_decoded_decoded_hi_lo_131 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_9_132 , core_csr_decoded_decoded_andMatrixInput_10_131 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_132 ={ core_csr_decoded_decoded_lo_lo_hi_125 , core_csr_decoded_decoded_andMatrixInput_11_125 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_132 ={ core_csr_decoded_decoded_andMatrixInput_6_132 , core_csr_decoded_decoded_andMatrixInput_7_132 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_133 ={ core_csr_decoded_decoded_lo_hi_hi_132 , core_csr_decoded_decoded_andMatrixInput_8_132 }; 
    wire[5:0] core_csr_decoded_decoded_lo_133 ={ core_csr_decoded_decoded_lo_hi_133 , core_csr_decoded_decoded_lo_lo_132 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_131 ={ core_csr_decoded_decoded_andMatrixInput_3_133 , core_csr_decoded_decoded_andMatrixInput_4_133 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_132 ={ core_csr_decoded_decoded_hi_lo_hi_131 , core_csr_decoded_decoded_andMatrixInput_5_133 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_132 ={ core_csr_decoded_decoded_andMatrixInput_0_133 , core_csr_decoded_decoded_andMatrixInput_1_133 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_133 ={ core_csr_decoded_decoded_hi_hi_hi_132 , core_csr_decoded_decoded_andMatrixInput_2_133 }; 
    wire[5:0] core_csr_decoded_decoded_hi_133 ={ core_csr_decoded_decoded_hi_hi_133 , core_csr_decoded_decoded_hi_lo_132 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_9_133 , core_csr_decoded_decoded_andMatrixInput_10_132 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_133 ={ core_csr_decoded_decoded_lo_lo_hi_126 , core_csr_decoded_decoded_andMatrixInput_11_126 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_133 ={ core_csr_decoded_decoded_andMatrixInput_6_133 , core_csr_decoded_decoded_andMatrixInput_7_133 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_134 ={ core_csr_decoded_decoded_lo_hi_hi_133 , core_csr_decoded_decoded_andMatrixInput_8_133 }; 
    wire[5:0] core_csr_decoded_decoded_lo_134 ={ core_csr_decoded_decoded_lo_hi_134 , core_csr_decoded_decoded_lo_lo_133 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_132 ={ core_csr_decoded_decoded_andMatrixInput_3_134 , core_csr_decoded_decoded_andMatrixInput_4_134 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_133 ={ core_csr_decoded_decoded_hi_lo_hi_132 , core_csr_decoded_decoded_andMatrixInput_5_134 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_133 ={ core_csr_decoded_decoded_andMatrixInput_0_134 , core_csr_decoded_decoded_andMatrixInput_1_134 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_134 ={ core_csr_decoded_decoded_hi_hi_hi_133 , core_csr_decoded_decoded_andMatrixInput_2_134 }; 
    wire[5:0] core_csr_decoded_decoded_hi_134 ={ core_csr_decoded_decoded_hi_hi_134 , core_csr_decoded_decoded_hi_lo_133 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_9_134 , core_csr_decoded_decoded_andMatrixInput_10_133 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_134 ={ core_csr_decoded_decoded_lo_lo_hi_127 , core_csr_decoded_decoded_andMatrixInput_11_127 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_134 ={ core_csr_decoded_decoded_andMatrixInput_6_134 , core_csr_decoded_decoded_andMatrixInput_7_134 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_135 ={ core_csr_decoded_decoded_lo_hi_hi_134 , core_csr_decoded_decoded_andMatrixInput_8_134 }; 
    wire[5:0] core_csr_decoded_decoded_lo_135 ={ core_csr_decoded_decoded_lo_hi_135 , core_csr_decoded_decoded_lo_lo_134 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_133 ={ core_csr_decoded_decoded_andMatrixInput_3_135 , core_csr_decoded_decoded_andMatrixInput_4_135 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_134 ={ core_csr_decoded_decoded_hi_lo_hi_133 , core_csr_decoded_decoded_andMatrixInput_5_135 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_134 ={ core_csr_decoded_decoded_andMatrixInput_0_135 , core_csr_decoded_decoded_andMatrixInput_1_135 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_135 ={ core_csr_decoded_decoded_hi_hi_hi_134 , core_csr_decoded_decoded_andMatrixInput_2_135 }; 
    wire[5:0] core_csr_decoded_decoded_hi_135 ={ core_csr_decoded_decoded_hi_hi_135 , core_csr_decoded_decoded_hi_lo_134 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_9_135 , core_csr_decoded_decoded_andMatrixInput_10_134 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_135 ={ core_csr_decoded_decoded_lo_lo_hi_128 , core_csr_decoded_decoded_andMatrixInput_11_128 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_135 ={ core_csr_decoded_decoded_andMatrixInput_6_135 , core_csr_decoded_decoded_andMatrixInput_7_135 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_136 ={ core_csr_decoded_decoded_lo_hi_hi_135 , core_csr_decoded_decoded_andMatrixInput_8_135 }; 
    wire[5:0] core_csr_decoded_decoded_lo_136 ={ core_csr_decoded_decoded_lo_hi_136 , core_csr_decoded_decoded_lo_lo_135 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_134 ={ core_csr_decoded_decoded_andMatrixInput_3_136 , core_csr_decoded_decoded_andMatrixInput_4_136 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_135 ={ core_csr_decoded_decoded_hi_lo_hi_134 , core_csr_decoded_decoded_andMatrixInput_5_136 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_135 ={ core_csr_decoded_decoded_andMatrixInput_0_136 , core_csr_decoded_decoded_andMatrixInput_1_136 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_136 ={ core_csr_decoded_decoded_hi_hi_hi_135 , core_csr_decoded_decoded_andMatrixInput_2_136 }; 
    wire[5:0] core_csr_decoded_decoded_hi_136 ={ core_csr_decoded_decoded_hi_hi_136 , core_csr_decoded_decoded_hi_lo_135 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_9_136 , core_csr_decoded_decoded_andMatrixInput_10_135 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_136 ={ core_csr_decoded_decoded_lo_lo_hi_129 , core_csr_decoded_decoded_andMatrixInput_11_129 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_136 ={ core_csr_decoded_decoded_andMatrixInput_6_136 , core_csr_decoded_decoded_andMatrixInput_7_136 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_137 ={ core_csr_decoded_decoded_lo_hi_hi_136 , core_csr_decoded_decoded_andMatrixInput_8_136 }; 
    wire[5:0] core_csr_decoded_decoded_lo_137 ={ core_csr_decoded_decoded_lo_hi_137 , core_csr_decoded_decoded_lo_lo_136 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_135 ={ core_csr_decoded_decoded_andMatrixInput_3_137 , core_csr_decoded_decoded_andMatrixInput_4_137 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_136 ={ core_csr_decoded_decoded_hi_lo_hi_135 , core_csr_decoded_decoded_andMatrixInput_5_137 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_136 ={ core_csr_decoded_decoded_andMatrixInput_0_137 , core_csr_decoded_decoded_andMatrixInput_1_137 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_137 ={ core_csr_decoded_decoded_hi_hi_hi_136 , core_csr_decoded_decoded_andMatrixInput_2_137 }; 
    wire[5:0] core_csr_decoded_decoded_hi_137 ={ core_csr_decoded_decoded_hi_hi_137 , core_csr_decoded_decoded_hi_lo_136 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_130 ={ core_csr_decoded_decoded_andMatrixInput_9_137 , core_csr_decoded_decoded_andMatrixInput_10_136 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_137 ={ core_csr_decoded_decoded_lo_lo_hi_130 , core_csr_decoded_decoded_andMatrixInput_11_130 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_137 ={ core_csr_decoded_decoded_andMatrixInput_6_137 , core_csr_decoded_decoded_andMatrixInput_7_137 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_138 ={ core_csr_decoded_decoded_lo_hi_hi_137 , core_csr_decoded_decoded_andMatrixInput_8_137 }; 
    wire[5:0] core_csr_decoded_decoded_lo_138 ={ core_csr_decoded_decoded_lo_hi_138 , core_csr_decoded_decoded_lo_lo_137 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_136 ={ core_csr_decoded_decoded_andMatrixInput_3_138 , core_csr_decoded_decoded_andMatrixInput_4_138 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_137 ={ core_csr_decoded_decoded_hi_lo_hi_136 , core_csr_decoded_decoded_andMatrixInput_5_138 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_137 ={ core_csr_decoded_decoded_andMatrixInput_0_138 , core_csr_decoded_decoded_andMatrixInput_1_138 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_138 ={ core_csr_decoded_decoded_hi_hi_hi_137 , core_csr_decoded_decoded_andMatrixInput_2_138 }; 
    wire[5:0] core_csr_decoded_decoded_hi_138 ={ core_csr_decoded_decoded_hi_hi_138 , core_csr_decoded_decoded_hi_lo_137 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_131 ={ core_csr_decoded_decoded_andMatrixInput_9_138 , core_csr_decoded_decoded_andMatrixInput_10_137 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_138 ={ core_csr_decoded_decoded_lo_lo_hi_131 , core_csr_decoded_decoded_andMatrixInput_11_131 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_138 ={ core_csr_decoded_decoded_andMatrixInput_6_138 , core_csr_decoded_decoded_andMatrixInput_7_138 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_139 ={ core_csr_decoded_decoded_lo_hi_hi_138 , core_csr_decoded_decoded_andMatrixInput_8_138 }; 
    wire[5:0] core_csr_decoded_decoded_lo_139 ={ core_csr_decoded_decoded_lo_hi_139 , core_csr_decoded_decoded_lo_lo_138 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_137 ={ core_csr_decoded_decoded_andMatrixInput_3_139 , core_csr_decoded_decoded_andMatrixInput_4_139 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_138 ={ core_csr_decoded_decoded_hi_lo_hi_137 , core_csr_decoded_decoded_andMatrixInput_5_139 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_138 ={ core_csr_decoded_decoded_andMatrixInput_0_139 , core_csr_decoded_decoded_andMatrixInput_1_139 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_139 ={ core_csr_decoded_decoded_hi_hi_hi_138 , core_csr_decoded_decoded_andMatrixInput_2_139 }; 
    wire[5:0] core_csr_decoded_decoded_hi_139 ={ core_csr_decoded_decoded_hi_hi_139 , core_csr_decoded_decoded_hi_lo_138 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_132 ={ core_csr_decoded_decoded_andMatrixInput_9_139 , core_csr_decoded_decoded_andMatrixInput_10_138 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_139 ={ core_csr_decoded_decoded_lo_lo_hi_132 , core_csr_decoded_decoded_andMatrixInput_11_132 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_139 ={ core_csr_decoded_decoded_andMatrixInput_6_139 , core_csr_decoded_decoded_andMatrixInput_7_139 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_140 ={ core_csr_decoded_decoded_lo_hi_hi_139 , core_csr_decoded_decoded_andMatrixInput_8_139 }; 
    wire[5:0] core_csr_decoded_decoded_lo_140 ={ core_csr_decoded_decoded_lo_hi_140 , core_csr_decoded_decoded_lo_lo_139 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_138 ={ core_csr_decoded_decoded_andMatrixInput_3_140 , core_csr_decoded_decoded_andMatrixInput_4_140 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_139 ={ core_csr_decoded_decoded_hi_lo_hi_138 , core_csr_decoded_decoded_andMatrixInput_5_140 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_139 ={ core_csr_decoded_decoded_andMatrixInput_0_140 , core_csr_decoded_decoded_andMatrixInput_1_140 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_140 ={ core_csr_decoded_decoded_hi_hi_hi_139 , core_csr_decoded_decoded_andMatrixInput_2_140 }; 
    wire[5:0] core_csr_decoded_decoded_hi_140 ={ core_csr_decoded_decoded_hi_hi_140 , core_csr_decoded_decoded_hi_lo_139 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_133 ={ core_csr_decoded_decoded_andMatrixInput_9_140 , core_csr_decoded_decoded_andMatrixInput_10_139 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_140 ={ core_csr_decoded_decoded_lo_lo_hi_133 , core_csr_decoded_decoded_andMatrixInput_11_133 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_140 ={ core_csr_decoded_decoded_andMatrixInput_6_140 , core_csr_decoded_decoded_andMatrixInput_7_140 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_141 ={ core_csr_decoded_decoded_lo_hi_hi_140 , core_csr_decoded_decoded_andMatrixInput_8_140 }; 
    wire[5:0] core_csr_decoded_decoded_lo_141 ={ core_csr_decoded_decoded_lo_hi_141 , core_csr_decoded_decoded_lo_lo_140 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_139 ={ core_csr_decoded_decoded_andMatrixInput_3_141 , core_csr_decoded_decoded_andMatrixInput_4_141 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_140 ={ core_csr_decoded_decoded_hi_lo_hi_139 , core_csr_decoded_decoded_andMatrixInput_5_141 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_140 ={ core_csr_decoded_decoded_andMatrixInput_0_141 , core_csr_decoded_decoded_andMatrixInput_1_141 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_141 ={ core_csr_decoded_decoded_hi_hi_hi_140 , core_csr_decoded_decoded_andMatrixInput_2_141 }; 
    wire[5:0] core_csr_decoded_decoded_hi_141 ={ core_csr_decoded_decoded_hi_hi_141 , core_csr_decoded_decoded_hi_lo_140 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_134 ={ core_csr_decoded_decoded_andMatrixInput_9_141 , core_csr_decoded_decoded_andMatrixInput_10_140 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_141 ={ core_csr_decoded_decoded_lo_lo_hi_134 , core_csr_decoded_decoded_andMatrixInput_11_134 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_141 ={ core_csr_decoded_decoded_andMatrixInput_6_141 , core_csr_decoded_decoded_andMatrixInput_7_141 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_142 ={ core_csr_decoded_decoded_lo_hi_hi_141 , core_csr_decoded_decoded_andMatrixInput_8_141 }; 
    wire[5:0] core_csr_decoded_decoded_lo_142 ={ core_csr_decoded_decoded_lo_hi_142 , core_csr_decoded_decoded_lo_lo_141 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_140 ={ core_csr_decoded_decoded_andMatrixInput_3_142 , core_csr_decoded_decoded_andMatrixInput_4_142 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_141 ={ core_csr_decoded_decoded_hi_lo_hi_140 , core_csr_decoded_decoded_andMatrixInput_5_142 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_141 ={ core_csr_decoded_decoded_andMatrixInput_0_142 , core_csr_decoded_decoded_andMatrixInput_1_142 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_142 ={ core_csr_decoded_decoded_hi_hi_hi_141 , core_csr_decoded_decoded_andMatrixInput_2_142 }; 
    wire[5:0] core_csr_decoded_decoded_hi_142 ={ core_csr_decoded_decoded_hi_hi_142 , core_csr_decoded_decoded_hi_lo_141 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_135 ={ core_csr_decoded_decoded_andMatrixInput_9_142 , core_csr_decoded_decoded_andMatrixInput_10_141 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_142 ={ core_csr_decoded_decoded_lo_lo_hi_135 , core_csr_decoded_decoded_andMatrixInput_11_135 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_142 ={ core_csr_decoded_decoded_andMatrixInput_6_142 , core_csr_decoded_decoded_andMatrixInput_7_142 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_143 ={ core_csr_decoded_decoded_lo_hi_hi_142 , core_csr_decoded_decoded_andMatrixInput_8_142 }; 
    wire[5:0] core_csr_decoded_decoded_lo_143 ={ core_csr_decoded_decoded_lo_hi_143 , core_csr_decoded_decoded_lo_lo_142 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_141 ={ core_csr_decoded_decoded_andMatrixInput_3_143 , core_csr_decoded_decoded_andMatrixInput_4_143 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_142 ={ core_csr_decoded_decoded_hi_lo_hi_141 , core_csr_decoded_decoded_andMatrixInput_5_143 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_142 ={ core_csr_decoded_decoded_andMatrixInput_0_143 , core_csr_decoded_decoded_andMatrixInput_1_143 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_143 ={ core_csr_decoded_decoded_hi_hi_hi_142 , core_csr_decoded_decoded_andMatrixInput_2_143 }; 
    wire[5:0] core_csr_decoded_decoded_hi_143 ={ core_csr_decoded_decoded_hi_hi_143 , core_csr_decoded_decoded_hi_lo_142 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_136 ={ core_csr_decoded_decoded_andMatrixInput_9_143 , core_csr_decoded_decoded_andMatrixInput_10_142 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_143 ={ core_csr_decoded_decoded_lo_lo_hi_136 , core_csr_decoded_decoded_andMatrixInput_11_136 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_143 ={ core_csr_decoded_decoded_andMatrixInput_6_143 , core_csr_decoded_decoded_andMatrixInput_7_143 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_144 ={ core_csr_decoded_decoded_lo_hi_hi_143 , core_csr_decoded_decoded_andMatrixInput_8_143 }; 
    wire[5:0] core_csr_decoded_decoded_lo_144 ={ core_csr_decoded_decoded_lo_hi_144 , core_csr_decoded_decoded_lo_lo_143 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_142 ={ core_csr_decoded_decoded_andMatrixInput_3_144 , core_csr_decoded_decoded_andMatrixInput_4_144 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_143 ={ core_csr_decoded_decoded_hi_lo_hi_142 , core_csr_decoded_decoded_andMatrixInput_5_144 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_143 ={ core_csr_decoded_decoded_andMatrixInput_0_144 , core_csr_decoded_decoded_andMatrixInput_1_144 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_144 ={ core_csr_decoded_decoded_hi_hi_hi_143 , core_csr_decoded_decoded_andMatrixInput_2_144 }; 
    wire[5:0] core_csr_decoded_decoded_hi_144 ={ core_csr_decoded_decoded_hi_hi_144 , core_csr_decoded_decoded_hi_lo_143 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_137 ={ core_csr_decoded_decoded_andMatrixInput_9_144 , core_csr_decoded_decoded_andMatrixInput_10_143 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_144 ={ core_csr_decoded_decoded_lo_lo_hi_137 , core_csr_decoded_decoded_andMatrixInput_11_137 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_144 ={ core_csr_decoded_decoded_andMatrixInput_6_144 , core_csr_decoded_decoded_andMatrixInput_7_144 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_145 ={ core_csr_decoded_decoded_lo_hi_hi_144 , core_csr_decoded_decoded_andMatrixInput_8_144 }; 
    wire[5:0] core_csr_decoded_decoded_lo_145 ={ core_csr_decoded_decoded_lo_hi_145 , core_csr_decoded_decoded_lo_lo_144 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_143 ={ core_csr_decoded_decoded_andMatrixInput_3_145 , core_csr_decoded_decoded_andMatrixInput_4_145 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_144 ={ core_csr_decoded_decoded_hi_lo_hi_143 , core_csr_decoded_decoded_andMatrixInput_5_145 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_144 ={ core_csr_decoded_decoded_andMatrixInput_0_145 , core_csr_decoded_decoded_andMatrixInput_1_145 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_145 ={ core_csr_decoded_decoded_hi_hi_hi_144 , core_csr_decoded_decoded_andMatrixInput_2_145 }; 
    wire[5:0] core_csr_decoded_decoded_hi_145 ={ core_csr_decoded_decoded_hi_hi_145 , core_csr_decoded_decoded_hi_lo_144 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_138 ={ core_csr_decoded_decoded_andMatrixInput_9_145 , core_csr_decoded_decoded_andMatrixInput_10_144 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_145 ={ core_csr_decoded_decoded_lo_lo_hi_138 , core_csr_decoded_decoded_andMatrixInput_11_138 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_145 ={ core_csr_decoded_decoded_andMatrixInput_6_145 , core_csr_decoded_decoded_andMatrixInput_7_145 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_146 ={ core_csr_decoded_decoded_lo_hi_hi_145 , core_csr_decoded_decoded_andMatrixInput_8_145 }; 
    wire[5:0] core_csr_decoded_decoded_lo_146 ={ core_csr_decoded_decoded_lo_hi_146 , core_csr_decoded_decoded_lo_lo_145 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_144 ={ core_csr_decoded_decoded_andMatrixInput_3_146 , core_csr_decoded_decoded_andMatrixInput_4_146 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_145 ={ core_csr_decoded_decoded_hi_lo_hi_144 , core_csr_decoded_decoded_andMatrixInput_5_146 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_145 ={ core_csr_decoded_decoded_andMatrixInput_0_146 , core_csr_decoded_decoded_andMatrixInput_1_146 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_146 ={ core_csr_decoded_decoded_hi_hi_hi_145 , core_csr_decoded_decoded_andMatrixInput_2_146 }; 
    wire[5:0] core_csr_decoded_decoded_hi_146 ={ core_csr_decoded_decoded_hi_hi_146 , core_csr_decoded_decoded_hi_lo_145 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_139 ={ core_csr_decoded_decoded_andMatrixInput_9_146 , core_csr_decoded_decoded_andMatrixInput_10_145 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_146 ={ core_csr_decoded_decoded_lo_lo_hi_139 , core_csr_decoded_decoded_andMatrixInput_11_139 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_146 ={ core_csr_decoded_decoded_andMatrixInput_6_146 , core_csr_decoded_decoded_andMatrixInput_7_146 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_147 ={ core_csr_decoded_decoded_lo_hi_hi_146 , core_csr_decoded_decoded_andMatrixInput_8_146 }; 
    wire[5:0] core_csr_decoded_decoded_lo_147 ={ core_csr_decoded_decoded_lo_hi_147 , core_csr_decoded_decoded_lo_lo_146 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_145 ={ core_csr_decoded_decoded_andMatrixInput_3_147 , core_csr_decoded_decoded_andMatrixInput_4_147 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_146 ={ core_csr_decoded_decoded_hi_lo_hi_145 , core_csr_decoded_decoded_andMatrixInput_5_147 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_146 ={ core_csr_decoded_decoded_andMatrixInput_0_147 , core_csr_decoded_decoded_andMatrixInput_1_147 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_147 ={ core_csr_decoded_decoded_hi_hi_hi_146 , core_csr_decoded_decoded_andMatrixInput_2_147 }; 
    wire[5:0] core_csr_decoded_decoded_hi_147 ={ core_csr_decoded_decoded_hi_hi_147 , core_csr_decoded_decoded_hi_lo_146 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_140 ={ core_csr_decoded_decoded_andMatrixInput_9_147 , core_csr_decoded_decoded_andMatrixInput_10_146 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_147 ={ core_csr_decoded_decoded_lo_lo_hi_140 , core_csr_decoded_decoded_andMatrixInput_11_140 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_147 ={ core_csr_decoded_decoded_andMatrixInput_6_147 , core_csr_decoded_decoded_andMatrixInput_7_147 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_148 ={ core_csr_decoded_decoded_lo_hi_hi_147 , core_csr_decoded_decoded_andMatrixInput_8_147 }; 
    wire[5:0] core_csr_decoded_decoded_lo_148 ={ core_csr_decoded_decoded_lo_hi_148 , core_csr_decoded_decoded_lo_lo_147 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_146 ={ core_csr_decoded_decoded_andMatrixInput_3_148 , core_csr_decoded_decoded_andMatrixInput_4_148 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_147 ={ core_csr_decoded_decoded_hi_lo_hi_146 , core_csr_decoded_decoded_andMatrixInput_5_148 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_147 ={ core_csr_decoded_decoded_andMatrixInput_0_148 , core_csr_decoded_decoded_andMatrixInput_1_148 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_148 ={ core_csr_decoded_decoded_hi_hi_hi_147 , core_csr_decoded_decoded_andMatrixInput_2_148 }; 
    wire[5:0] core_csr_decoded_decoded_hi_148 ={ core_csr_decoded_decoded_hi_hi_148 , core_csr_decoded_decoded_hi_lo_147 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_141 ={ core_csr_decoded_decoded_andMatrixInput_9_148 , core_csr_decoded_decoded_andMatrixInput_10_147 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_148 ={ core_csr_decoded_decoded_lo_lo_hi_141 , core_csr_decoded_decoded_andMatrixInput_11_141 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_148 ={ core_csr_decoded_decoded_andMatrixInput_6_148 , core_csr_decoded_decoded_andMatrixInput_7_148 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_149 ={ core_csr_decoded_decoded_lo_hi_hi_148 , core_csr_decoded_decoded_andMatrixInput_8_148 }; 
    wire[5:0] core_csr_decoded_decoded_lo_149 ={ core_csr_decoded_decoded_lo_hi_149 , core_csr_decoded_decoded_lo_lo_148 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_147 ={ core_csr_decoded_decoded_andMatrixInput_3_149 , core_csr_decoded_decoded_andMatrixInput_4_149 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_148 ={ core_csr_decoded_decoded_hi_lo_hi_147 , core_csr_decoded_decoded_andMatrixInput_5_149 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_148 ={ core_csr_decoded_decoded_andMatrixInput_0_149 , core_csr_decoded_decoded_andMatrixInput_1_149 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_149 ={ core_csr_decoded_decoded_hi_hi_hi_148 , core_csr_decoded_decoded_andMatrixInput_2_149 }; 
    wire[5:0] core_csr_decoded_decoded_hi_149 ={ core_csr_decoded_decoded_hi_hi_149 , core_csr_decoded_decoded_hi_lo_148 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_142 ={ core_csr_decoded_decoded_andMatrixInput_9_149 , core_csr_decoded_decoded_andMatrixInput_10_148 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_149 ={ core_csr_decoded_decoded_lo_lo_hi_142 , core_csr_decoded_decoded_andMatrixInput_11_142 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_149 ={ core_csr_decoded_decoded_andMatrixInput_6_149 , core_csr_decoded_decoded_andMatrixInput_7_149 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_150 ={ core_csr_decoded_decoded_lo_hi_hi_149 , core_csr_decoded_decoded_andMatrixInput_8_149 }; 
    wire[5:0] core_csr_decoded_decoded_lo_150 ={ core_csr_decoded_decoded_lo_hi_150 , core_csr_decoded_decoded_lo_lo_149 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_148 ={ core_csr_decoded_decoded_andMatrixInput_3_150 , core_csr_decoded_decoded_andMatrixInput_4_150 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_149 ={ core_csr_decoded_decoded_hi_lo_hi_148 , core_csr_decoded_decoded_andMatrixInput_5_150 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_149 ={ core_csr_decoded_decoded_andMatrixInput_0_150 , core_csr_decoded_decoded_andMatrixInput_1_150 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_150 ={ core_csr_decoded_decoded_hi_hi_hi_149 , core_csr_decoded_decoded_andMatrixInput_2_150 }; 
    wire[5:0] core_csr_decoded_decoded_hi_150 ={ core_csr_decoded_decoded_hi_hi_150 , core_csr_decoded_decoded_hi_lo_149 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_143 ={ core_csr_decoded_decoded_andMatrixInput_9_150 , core_csr_decoded_decoded_andMatrixInput_10_149 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_150 ={ core_csr_decoded_decoded_lo_lo_hi_143 , core_csr_decoded_decoded_andMatrixInput_11_143 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_150 ={ core_csr_decoded_decoded_andMatrixInput_6_150 , core_csr_decoded_decoded_andMatrixInput_7_150 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_151 ={ core_csr_decoded_decoded_lo_hi_hi_150 , core_csr_decoded_decoded_andMatrixInput_8_150 }; 
    wire[5:0] core_csr_decoded_decoded_lo_151 ={ core_csr_decoded_decoded_lo_hi_151 , core_csr_decoded_decoded_lo_lo_150 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_149 ={ core_csr_decoded_decoded_andMatrixInput_3_151 , core_csr_decoded_decoded_andMatrixInput_4_151 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_150 ={ core_csr_decoded_decoded_hi_lo_hi_149 , core_csr_decoded_decoded_andMatrixInput_5_151 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_150 ={ core_csr_decoded_decoded_andMatrixInput_0_151 , core_csr_decoded_decoded_andMatrixInput_1_151 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_151 ={ core_csr_decoded_decoded_hi_hi_hi_150 , core_csr_decoded_decoded_andMatrixInput_2_151 }; 
    wire[5:0] core_csr_decoded_decoded_hi_151 ={ core_csr_decoded_decoded_hi_hi_151 , core_csr_decoded_decoded_hi_lo_150 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_144 ={ core_csr_decoded_decoded_andMatrixInput_9_151 , core_csr_decoded_decoded_andMatrixInput_10_150 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_151 ={ core_csr_decoded_decoded_lo_lo_hi_144 , core_csr_decoded_decoded_andMatrixInput_11_144 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_151 ={ core_csr_decoded_decoded_andMatrixInput_6_151 , core_csr_decoded_decoded_andMatrixInput_7_151 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_152 ={ core_csr_decoded_decoded_lo_hi_hi_151 , core_csr_decoded_decoded_andMatrixInput_8_151 }; 
    wire[5:0] core_csr_decoded_decoded_lo_152 ={ core_csr_decoded_decoded_lo_hi_152 , core_csr_decoded_decoded_lo_lo_151 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_150 ={ core_csr_decoded_decoded_andMatrixInput_3_152 , core_csr_decoded_decoded_andMatrixInput_4_152 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_151 ={ core_csr_decoded_decoded_hi_lo_hi_150 , core_csr_decoded_decoded_andMatrixInput_5_152 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_151 ={ core_csr_decoded_decoded_andMatrixInput_0_152 , core_csr_decoded_decoded_andMatrixInput_1_152 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_152 ={ core_csr_decoded_decoded_hi_hi_hi_151 , core_csr_decoded_decoded_andMatrixInput_2_152 }; 
    wire[5:0] core_csr_decoded_decoded_hi_152 ={ core_csr_decoded_decoded_hi_hi_152 , core_csr_decoded_decoded_hi_lo_151 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_145 ={ core_csr_decoded_decoded_andMatrixInput_9_152 , core_csr_decoded_decoded_andMatrixInput_10_151 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_152 ={ core_csr_decoded_decoded_lo_lo_hi_145 , core_csr_decoded_decoded_andMatrixInput_11_145 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_152 ={ core_csr_decoded_decoded_andMatrixInput_6_152 , core_csr_decoded_decoded_andMatrixInput_7_152 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_153 ={ core_csr_decoded_decoded_lo_hi_hi_152 , core_csr_decoded_decoded_andMatrixInput_8_152 }; 
    wire[5:0] core_csr_decoded_decoded_lo_153 ={ core_csr_decoded_decoded_lo_hi_153 , core_csr_decoded_decoded_lo_lo_152 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_151 ={ core_csr_decoded_decoded_andMatrixInput_3_153 , core_csr_decoded_decoded_andMatrixInput_4_153 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_152 ={ core_csr_decoded_decoded_hi_lo_hi_151 , core_csr_decoded_decoded_andMatrixInput_5_153 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_152 ={ core_csr_decoded_decoded_andMatrixInput_0_153 , core_csr_decoded_decoded_andMatrixInput_1_153 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_153 ={ core_csr_decoded_decoded_hi_hi_hi_152 , core_csr_decoded_decoded_andMatrixInput_2_153 }; 
    wire[5:0] core_csr_decoded_decoded_hi_153 ={ core_csr_decoded_decoded_hi_hi_153 , core_csr_decoded_decoded_hi_lo_152 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_146 ={ core_csr_decoded_decoded_andMatrixInput_9_153 , core_csr_decoded_decoded_andMatrixInput_10_152 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_153 ={ core_csr_decoded_decoded_lo_lo_hi_146 , core_csr_decoded_decoded_andMatrixInput_11_146 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_153 ={ core_csr_decoded_decoded_andMatrixInput_6_153 , core_csr_decoded_decoded_andMatrixInput_7_153 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_154 ={ core_csr_decoded_decoded_lo_hi_hi_153 , core_csr_decoded_decoded_andMatrixInput_8_153 }; 
    wire[5:0] core_csr_decoded_decoded_lo_154 ={ core_csr_decoded_decoded_lo_hi_154 , core_csr_decoded_decoded_lo_lo_153 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_152 ={ core_csr_decoded_decoded_andMatrixInput_3_154 , core_csr_decoded_decoded_andMatrixInput_4_154 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_153 ={ core_csr_decoded_decoded_hi_lo_hi_152 , core_csr_decoded_decoded_andMatrixInput_5_154 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_153 ={ core_csr_decoded_decoded_andMatrixInput_0_154 , core_csr_decoded_decoded_andMatrixInput_1_154 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_154 ={ core_csr_decoded_decoded_hi_hi_hi_153 , core_csr_decoded_decoded_andMatrixInput_2_154 }; 
    wire[5:0] core_csr_decoded_decoded_hi_154 ={ core_csr_decoded_decoded_hi_hi_154 , core_csr_decoded_decoded_hi_lo_153 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_147 ={ core_csr_decoded_decoded_andMatrixInput_9_154 , core_csr_decoded_decoded_andMatrixInput_10_153 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_154 ={ core_csr_decoded_decoded_lo_lo_hi_147 , core_csr_decoded_decoded_andMatrixInput_11_147 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_154 ={ core_csr_decoded_decoded_andMatrixInput_6_154 , core_csr_decoded_decoded_andMatrixInput_7_154 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_155 ={ core_csr_decoded_decoded_lo_hi_hi_154 , core_csr_decoded_decoded_andMatrixInput_8_154 }; 
    wire[5:0] core_csr_decoded_decoded_lo_155 ={ core_csr_decoded_decoded_lo_hi_155 , core_csr_decoded_decoded_lo_lo_154 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_153 ={ core_csr_decoded_decoded_andMatrixInput_3_155 , core_csr_decoded_decoded_andMatrixInput_4_155 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_154 ={ core_csr_decoded_decoded_hi_lo_hi_153 , core_csr_decoded_decoded_andMatrixInput_5_155 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_154 ={ core_csr_decoded_decoded_andMatrixInput_0_155 , core_csr_decoded_decoded_andMatrixInput_1_155 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_155 ={ core_csr_decoded_decoded_hi_hi_hi_154 , core_csr_decoded_decoded_andMatrixInput_2_155 }; 
    wire[5:0] core_csr_decoded_decoded_hi_155 ={ core_csr_decoded_decoded_hi_hi_155 , core_csr_decoded_decoded_hi_lo_154 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_148 ={ core_csr_decoded_decoded_andMatrixInput_9_155 , core_csr_decoded_decoded_andMatrixInput_10_154 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_155 ={ core_csr_decoded_decoded_lo_lo_hi_148 , core_csr_decoded_decoded_andMatrixInput_11_148 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_155 ={ core_csr_decoded_decoded_andMatrixInput_6_155 , core_csr_decoded_decoded_andMatrixInput_7_155 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_156 ={ core_csr_decoded_decoded_lo_hi_hi_155 , core_csr_decoded_decoded_andMatrixInput_8_155 }; 
    wire[5:0] core_csr_decoded_decoded_lo_156 ={ core_csr_decoded_decoded_lo_hi_156 , core_csr_decoded_decoded_lo_lo_155 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_154 ={ core_csr_decoded_decoded_andMatrixInput_3_156 , core_csr_decoded_decoded_andMatrixInput_4_156 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_155 ={ core_csr_decoded_decoded_hi_lo_hi_154 , core_csr_decoded_decoded_andMatrixInput_5_156 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_155 ={ core_csr_decoded_decoded_andMatrixInput_0_156 , core_csr_decoded_decoded_andMatrixInput_1_156 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_156 ={ core_csr_decoded_decoded_hi_hi_hi_155 , core_csr_decoded_decoded_andMatrixInput_2_156 }; 
    wire[5:0] core_csr_decoded_decoded_hi_156 ={ core_csr_decoded_decoded_hi_hi_156 , core_csr_decoded_decoded_hi_lo_155 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_149 ={ core_csr_decoded_decoded_andMatrixInput_9_156 , core_csr_decoded_decoded_andMatrixInput_10_155 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_156 ={ core_csr_decoded_decoded_lo_lo_hi_149 , core_csr_decoded_decoded_andMatrixInput_11_149 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_156 ={ core_csr_decoded_decoded_andMatrixInput_6_156 , core_csr_decoded_decoded_andMatrixInput_7_156 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_157 ={ core_csr_decoded_decoded_lo_hi_hi_156 , core_csr_decoded_decoded_andMatrixInput_8_156 }; 
    wire[5:0] core_csr_decoded_decoded_lo_157 ={ core_csr_decoded_decoded_lo_hi_157 , core_csr_decoded_decoded_lo_lo_156 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_155 ={ core_csr_decoded_decoded_andMatrixInput_3_157 , core_csr_decoded_decoded_andMatrixInput_4_157 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_156 ={ core_csr_decoded_decoded_hi_lo_hi_155 , core_csr_decoded_decoded_andMatrixInput_5_157 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_156 ={ core_csr_decoded_decoded_andMatrixInput_0_157 , core_csr_decoded_decoded_andMatrixInput_1_157 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_157 ={ core_csr_decoded_decoded_hi_hi_hi_156 , core_csr_decoded_decoded_andMatrixInput_2_157 }; 
    wire[5:0] core_csr_decoded_decoded_hi_157 ={ core_csr_decoded_decoded_hi_hi_157 , core_csr_decoded_decoded_hi_lo_156 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_150 ={ core_csr_decoded_decoded_andMatrixInput_9_157 , core_csr_decoded_decoded_andMatrixInput_10_156 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_157 ={ core_csr_decoded_decoded_lo_lo_hi_150 , core_csr_decoded_decoded_andMatrixInput_11_150 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_157 ={ core_csr_decoded_decoded_andMatrixInput_6_157 , core_csr_decoded_decoded_andMatrixInput_7_157 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_158 ={ core_csr_decoded_decoded_lo_hi_hi_157 , core_csr_decoded_decoded_andMatrixInput_8_157 }; 
    wire[5:0] core_csr_decoded_decoded_lo_158 ={ core_csr_decoded_decoded_lo_hi_158 , core_csr_decoded_decoded_lo_lo_157 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_156 ={ core_csr_decoded_decoded_andMatrixInput_3_158 , core_csr_decoded_decoded_andMatrixInput_4_158 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_157 ={ core_csr_decoded_decoded_hi_lo_hi_156 , core_csr_decoded_decoded_andMatrixInput_5_158 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_157 ={ core_csr_decoded_decoded_andMatrixInput_0_158 , core_csr_decoded_decoded_andMatrixInput_1_158 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_158 ={ core_csr_decoded_decoded_hi_hi_hi_157 , core_csr_decoded_decoded_andMatrixInput_2_158 }; 
    wire[5:0] core_csr_decoded_decoded_hi_158 ={ core_csr_decoded_decoded_hi_hi_158 , core_csr_decoded_decoded_hi_lo_157 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_151 ={ core_csr_decoded_decoded_andMatrixInput_9_158 , core_csr_decoded_decoded_andMatrixInput_10_157 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_158 ={ core_csr_decoded_decoded_lo_lo_hi_151 , core_csr_decoded_decoded_andMatrixInput_11_151 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_158 ={ core_csr_decoded_decoded_andMatrixInput_6_158 , core_csr_decoded_decoded_andMatrixInput_7_158 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_159 ={ core_csr_decoded_decoded_lo_hi_hi_158 , core_csr_decoded_decoded_andMatrixInput_8_158 }; 
    wire[5:0] core_csr_decoded_decoded_lo_159 ={ core_csr_decoded_decoded_lo_hi_159 , core_csr_decoded_decoded_lo_lo_158 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_157 ={ core_csr_decoded_decoded_andMatrixInput_3_159 , core_csr_decoded_decoded_andMatrixInput_4_159 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_158 ={ core_csr_decoded_decoded_hi_lo_hi_157 , core_csr_decoded_decoded_andMatrixInput_5_159 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_158 ={ core_csr_decoded_decoded_andMatrixInput_0_159 , core_csr_decoded_decoded_andMatrixInput_1_159 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_159 ={ core_csr_decoded_decoded_hi_hi_hi_158 , core_csr_decoded_decoded_andMatrixInput_2_159 }; 
    wire[5:0] core_csr_decoded_decoded_hi_159 ={ core_csr_decoded_decoded_hi_hi_159 , core_csr_decoded_decoded_hi_lo_158 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_159 ={ core_csr_decoded_decoded_andMatrixInput_9_159 , core_csr_decoded_decoded_andMatrixInput_10_158 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_159 ={ core_csr_decoded_decoded_andMatrixInput_6_159 , core_csr_decoded_decoded_andMatrixInput_7_159 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_160 ={ core_csr_decoded_decoded_lo_hi_hi_159 , core_csr_decoded_decoded_andMatrixInput_8_159 }; 
    wire[4:0] core_csr_decoded_decoded_lo_160 ={ core_csr_decoded_decoded_lo_hi_160 , core_csr_decoded_decoded_lo_lo_159 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_158 ={ core_csr_decoded_decoded_andMatrixInput_3_160 , core_csr_decoded_decoded_andMatrixInput_4_160 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_159 ={ core_csr_decoded_decoded_hi_lo_hi_158 , core_csr_decoded_decoded_andMatrixInput_5_160 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_159 ={ core_csr_decoded_decoded_andMatrixInput_0_160 , core_csr_decoded_decoded_andMatrixInput_1_160 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_160 ={ core_csr_decoded_decoded_hi_hi_hi_159 , core_csr_decoded_decoded_andMatrixInput_2_160 }; 
    wire[5:0] core_csr_decoded_decoded_hi_160 ={ core_csr_decoded_decoded_hi_hi_160 , core_csr_decoded_decoded_hi_lo_159 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_152 ={ core_csr_decoded_decoded_andMatrixInput_9_160 , core_csr_decoded_decoded_andMatrixInput_10_159 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_160 ={ core_csr_decoded_decoded_lo_lo_hi_152 , core_csr_decoded_decoded_andMatrixInput_11_152 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_160 ={ core_csr_decoded_decoded_andMatrixInput_6_160 , core_csr_decoded_decoded_andMatrixInput_7_160 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_161 ={ core_csr_decoded_decoded_lo_hi_hi_160 , core_csr_decoded_decoded_andMatrixInput_8_160 }; 
    wire[5:0] core_csr_decoded_decoded_lo_161 ={ core_csr_decoded_decoded_lo_hi_161 , core_csr_decoded_decoded_lo_lo_160 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_159 ={ core_csr_decoded_decoded_andMatrixInput_3_161 , core_csr_decoded_decoded_andMatrixInput_4_161 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_160 ={ core_csr_decoded_decoded_hi_lo_hi_159 , core_csr_decoded_decoded_andMatrixInput_5_161 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_160 ={ core_csr_decoded_decoded_andMatrixInput_0_161 , core_csr_decoded_decoded_andMatrixInput_1_161 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_161 ={ core_csr_decoded_decoded_hi_hi_hi_160 , core_csr_decoded_decoded_andMatrixInput_2_161 }; 
    wire[5:0] core_csr_decoded_decoded_hi_161 ={ core_csr_decoded_decoded_hi_hi_161 , core_csr_decoded_decoded_hi_lo_160 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_153 ={ core_csr_decoded_decoded_andMatrixInput_9_161 , core_csr_decoded_decoded_andMatrixInput_10_160 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_161 ={ core_csr_decoded_decoded_lo_lo_hi_153 , core_csr_decoded_decoded_andMatrixInput_11_153 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_161 ={ core_csr_decoded_decoded_andMatrixInput_6_161 , core_csr_decoded_decoded_andMatrixInput_7_161 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_162 ={ core_csr_decoded_decoded_lo_hi_hi_161 , core_csr_decoded_decoded_andMatrixInput_8_161 }; 
    wire[5:0] core_csr_decoded_decoded_lo_162 ={ core_csr_decoded_decoded_lo_hi_162 , core_csr_decoded_decoded_lo_lo_161 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_160 ={ core_csr_decoded_decoded_andMatrixInput_3_162 , core_csr_decoded_decoded_andMatrixInput_4_162 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_161 ={ core_csr_decoded_decoded_hi_lo_hi_160 , core_csr_decoded_decoded_andMatrixInput_5_162 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_161 ={ core_csr_decoded_decoded_andMatrixInput_0_162 , core_csr_decoded_decoded_andMatrixInput_1_162 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_162 ={ core_csr_decoded_decoded_hi_hi_hi_161 , core_csr_decoded_decoded_andMatrixInput_2_162 }; 
    wire[5:0] core_csr_decoded_decoded_hi_162 ={ core_csr_decoded_decoded_hi_hi_162 , core_csr_decoded_decoded_hi_lo_161 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_154 ={ core_csr_decoded_decoded_andMatrixInput_9_162 , core_csr_decoded_decoded_andMatrixInput_10_161 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_162 ={ core_csr_decoded_decoded_lo_lo_hi_154 , core_csr_decoded_decoded_andMatrixInput_11_154 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_162 ={ core_csr_decoded_decoded_andMatrixInput_6_162 , core_csr_decoded_decoded_andMatrixInput_7_162 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_163 ={ core_csr_decoded_decoded_lo_hi_hi_162 , core_csr_decoded_decoded_andMatrixInput_8_162 }; 
    wire[5:0] core_csr_decoded_decoded_lo_163 ={ core_csr_decoded_decoded_lo_hi_163 , core_csr_decoded_decoded_lo_lo_162 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_161 ={ core_csr_decoded_decoded_andMatrixInput_3_163 , core_csr_decoded_decoded_andMatrixInput_4_163 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_162 ={ core_csr_decoded_decoded_hi_lo_hi_161 , core_csr_decoded_decoded_andMatrixInput_5_163 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_162 ={ core_csr_decoded_decoded_andMatrixInput_0_163 , core_csr_decoded_decoded_andMatrixInput_1_163 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_163 ={ core_csr_decoded_decoded_hi_hi_hi_162 , core_csr_decoded_decoded_andMatrixInput_2_163 }; 
    wire[5:0] core_csr_decoded_decoded_hi_163 ={ core_csr_decoded_decoded_hi_hi_163 , core_csr_decoded_decoded_hi_lo_162 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_155 ={ core_csr_decoded_decoded_andMatrixInput_9_163 , core_csr_decoded_decoded_andMatrixInput_10_162 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_163 ={ core_csr_decoded_decoded_lo_lo_hi_155 , core_csr_decoded_decoded_andMatrixInput_11_155 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_163 ={ core_csr_decoded_decoded_andMatrixInput_6_163 , core_csr_decoded_decoded_andMatrixInput_7_163 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_164 ={ core_csr_decoded_decoded_lo_hi_hi_163 , core_csr_decoded_decoded_andMatrixInput_8_163 }; 
    wire[5:0] core_csr_decoded_decoded_lo_164 ={ core_csr_decoded_decoded_lo_hi_164 , core_csr_decoded_decoded_lo_lo_163 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_162 ={ core_csr_decoded_decoded_andMatrixInput_3_164 , core_csr_decoded_decoded_andMatrixInput_4_164 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_163 ={ core_csr_decoded_decoded_hi_lo_hi_162 , core_csr_decoded_decoded_andMatrixInput_5_164 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_163 ={ core_csr_decoded_decoded_andMatrixInput_0_164 , core_csr_decoded_decoded_andMatrixInput_1_164 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_164 ={ core_csr_decoded_decoded_hi_hi_hi_163 , core_csr_decoded_decoded_andMatrixInput_2_164 }; 
    wire[5:0] core_csr_decoded_decoded_hi_164 ={ core_csr_decoded_decoded_hi_hi_164 , core_csr_decoded_decoded_hi_lo_163 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_156 ={ core_csr_decoded_decoded_andMatrixInput_9_164 , core_csr_decoded_decoded_andMatrixInput_10_163 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_164 ={ core_csr_decoded_decoded_lo_lo_hi_156 , core_csr_decoded_decoded_andMatrixInput_11_156 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_164 ={ core_csr_decoded_decoded_andMatrixInput_6_164 , core_csr_decoded_decoded_andMatrixInput_7_164 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_165 ={ core_csr_decoded_decoded_lo_hi_hi_164 , core_csr_decoded_decoded_andMatrixInput_8_164 }; 
    wire[5:0] core_csr_decoded_decoded_lo_165 ={ core_csr_decoded_decoded_lo_hi_165 , core_csr_decoded_decoded_lo_lo_164 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_163 ={ core_csr_decoded_decoded_andMatrixInput_3_165 , core_csr_decoded_decoded_andMatrixInput_4_165 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_164 ={ core_csr_decoded_decoded_hi_lo_hi_163 , core_csr_decoded_decoded_andMatrixInput_5_165 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_164 ={ core_csr_decoded_decoded_andMatrixInput_0_165 , core_csr_decoded_decoded_andMatrixInput_1_165 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_165 ={ core_csr_decoded_decoded_hi_hi_hi_164 , core_csr_decoded_decoded_andMatrixInput_2_165 }; 
    wire[5:0] core_csr_decoded_decoded_hi_165 ={ core_csr_decoded_decoded_hi_hi_165 , core_csr_decoded_decoded_hi_lo_164 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_157 ={ core_csr_decoded_decoded_andMatrixInput_9_165 , core_csr_decoded_decoded_andMatrixInput_10_164 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_165 ={ core_csr_decoded_decoded_lo_lo_hi_157 , core_csr_decoded_decoded_andMatrixInput_11_157 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_165 ={ core_csr_decoded_decoded_andMatrixInput_6_165 , core_csr_decoded_decoded_andMatrixInput_7_165 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_166 ={ core_csr_decoded_decoded_lo_hi_hi_165 , core_csr_decoded_decoded_andMatrixInput_8_165 }; 
    wire[5:0] core_csr_decoded_decoded_lo_166 ={ core_csr_decoded_decoded_lo_hi_166 , core_csr_decoded_decoded_lo_lo_165 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_164 ={ core_csr_decoded_decoded_andMatrixInput_3_166 , core_csr_decoded_decoded_andMatrixInput_4_166 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_165 ={ core_csr_decoded_decoded_hi_lo_hi_164 , core_csr_decoded_decoded_andMatrixInput_5_166 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_165 ={ core_csr_decoded_decoded_andMatrixInput_0_166 , core_csr_decoded_decoded_andMatrixInput_1_166 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_166 ={ core_csr_decoded_decoded_hi_hi_hi_165 , core_csr_decoded_decoded_andMatrixInput_2_166 }; 
    wire[5:0] core_csr_decoded_decoded_hi_166 ={ core_csr_decoded_decoded_hi_hi_166 , core_csr_decoded_decoded_hi_lo_165 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_158 ={ core_csr_decoded_decoded_andMatrixInput_9_166 , core_csr_decoded_decoded_andMatrixInput_10_165 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_166 ={ core_csr_decoded_decoded_lo_lo_hi_158 , core_csr_decoded_decoded_andMatrixInput_11_158 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_166 ={ core_csr_decoded_decoded_andMatrixInput_6_166 , core_csr_decoded_decoded_andMatrixInput_7_166 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_167 ={ core_csr_decoded_decoded_lo_hi_hi_166 , core_csr_decoded_decoded_andMatrixInput_8_166 }; 
    wire[5:0] core_csr_decoded_decoded_lo_167 ={ core_csr_decoded_decoded_lo_hi_167 , core_csr_decoded_decoded_lo_lo_166 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_165 ={ core_csr_decoded_decoded_andMatrixInput_3_167 , core_csr_decoded_decoded_andMatrixInput_4_167 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_166 ={ core_csr_decoded_decoded_hi_lo_hi_165 , core_csr_decoded_decoded_andMatrixInput_5_167 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_166 ={ core_csr_decoded_decoded_andMatrixInput_0_167 , core_csr_decoded_decoded_andMatrixInput_1_167 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_167 ={ core_csr_decoded_decoded_hi_hi_hi_166 , core_csr_decoded_decoded_andMatrixInput_2_167 }; 
    wire[5:0] core_csr_decoded_decoded_hi_167 ={ core_csr_decoded_decoded_hi_hi_167 , core_csr_decoded_decoded_hi_lo_166 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_159 ={ core_csr_decoded_decoded_andMatrixInput_9_167 , core_csr_decoded_decoded_andMatrixInput_10_166 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_167 ={ core_csr_decoded_decoded_lo_lo_hi_159 , core_csr_decoded_decoded_andMatrixInput_11_159 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_167 ={ core_csr_decoded_decoded_andMatrixInput_6_167 , core_csr_decoded_decoded_andMatrixInput_7_167 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_168 ={ core_csr_decoded_decoded_lo_hi_hi_167 , core_csr_decoded_decoded_andMatrixInput_8_167 }; 
    wire[5:0] core_csr_decoded_decoded_lo_168 ={ core_csr_decoded_decoded_lo_hi_168 , core_csr_decoded_decoded_lo_lo_167 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_166 ={ core_csr_decoded_decoded_andMatrixInput_3_168 , core_csr_decoded_decoded_andMatrixInput_4_168 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_167 ={ core_csr_decoded_decoded_hi_lo_hi_166 , core_csr_decoded_decoded_andMatrixInput_5_168 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_167 ={ core_csr_decoded_decoded_andMatrixInput_0_168 , core_csr_decoded_decoded_andMatrixInput_1_168 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_168 ={ core_csr_decoded_decoded_hi_hi_hi_167 , core_csr_decoded_decoded_andMatrixInput_2_168 }; 
    wire[5:0] core_csr_decoded_decoded_hi_168 ={ core_csr_decoded_decoded_hi_hi_168 , core_csr_decoded_decoded_hi_lo_167 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_160 ={ core_csr_decoded_decoded_andMatrixInput_9_168 , core_csr_decoded_decoded_andMatrixInput_10_167 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_168 ={ core_csr_decoded_decoded_lo_lo_hi_160 , core_csr_decoded_decoded_andMatrixInput_11_160 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_168 ={ core_csr_decoded_decoded_andMatrixInput_6_168 , core_csr_decoded_decoded_andMatrixInput_7_168 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_169 ={ core_csr_decoded_decoded_lo_hi_hi_168 , core_csr_decoded_decoded_andMatrixInput_8_168 }; 
    wire[5:0] core_csr_decoded_decoded_lo_169 ={ core_csr_decoded_decoded_lo_hi_169 , core_csr_decoded_decoded_lo_lo_168 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_167 ={ core_csr_decoded_decoded_andMatrixInput_3_169 , core_csr_decoded_decoded_andMatrixInput_4_169 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_168 ={ core_csr_decoded_decoded_hi_lo_hi_167 , core_csr_decoded_decoded_andMatrixInput_5_169 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_168 ={ core_csr_decoded_decoded_andMatrixInput_0_169 , core_csr_decoded_decoded_andMatrixInput_1_169 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_169 ={ core_csr_decoded_decoded_hi_hi_hi_168 , core_csr_decoded_decoded_andMatrixInput_2_169 }; 
    wire[5:0] core_csr_decoded_decoded_hi_169 ={ core_csr_decoded_decoded_hi_hi_169 , core_csr_decoded_decoded_hi_lo_168 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_161 ={ core_csr_decoded_decoded_andMatrixInput_9_169 , core_csr_decoded_decoded_andMatrixInput_10_168 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_169 ={ core_csr_decoded_decoded_lo_lo_hi_161 , core_csr_decoded_decoded_andMatrixInput_11_161 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_169 ={ core_csr_decoded_decoded_andMatrixInput_6_169 , core_csr_decoded_decoded_andMatrixInput_7_169 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_170 ={ core_csr_decoded_decoded_lo_hi_hi_169 , core_csr_decoded_decoded_andMatrixInput_8_169 }; 
    wire[5:0] core_csr_decoded_decoded_lo_170 ={ core_csr_decoded_decoded_lo_hi_170 , core_csr_decoded_decoded_lo_lo_169 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_168 ={ core_csr_decoded_decoded_andMatrixInput_3_170 , core_csr_decoded_decoded_andMatrixInput_4_170 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_169 ={ core_csr_decoded_decoded_hi_lo_hi_168 , core_csr_decoded_decoded_andMatrixInput_5_170 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_169 ={ core_csr_decoded_decoded_andMatrixInput_0_170 , core_csr_decoded_decoded_andMatrixInput_1_170 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_170 ={ core_csr_decoded_decoded_hi_hi_hi_169 , core_csr_decoded_decoded_andMatrixInput_2_170 }; 
    wire[5:0] core_csr_decoded_decoded_hi_170 ={ core_csr_decoded_decoded_hi_hi_170 , core_csr_decoded_decoded_hi_lo_169 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_162 ={ core_csr_decoded_decoded_andMatrixInput_9_170 , core_csr_decoded_decoded_andMatrixInput_10_169 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_170 ={ core_csr_decoded_decoded_lo_lo_hi_162 , core_csr_decoded_decoded_andMatrixInput_11_162 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_170 ={ core_csr_decoded_decoded_andMatrixInput_6_170 , core_csr_decoded_decoded_andMatrixInput_7_170 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_171 ={ core_csr_decoded_decoded_lo_hi_hi_170 , core_csr_decoded_decoded_andMatrixInput_8_170 }; 
    wire[5:0] core_csr_decoded_decoded_lo_171 ={ core_csr_decoded_decoded_lo_hi_171 , core_csr_decoded_decoded_lo_lo_170 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_169 ={ core_csr_decoded_decoded_andMatrixInput_3_171 , core_csr_decoded_decoded_andMatrixInput_4_171 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_170 ={ core_csr_decoded_decoded_hi_lo_hi_169 , core_csr_decoded_decoded_andMatrixInput_5_171 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_170 ={ core_csr_decoded_decoded_andMatrixInput_0_171 , core_csr_decoded_decoded_andMatrixInput_1_171 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_171 ={ core_csr_decoded_decoded_hi_hi_hi_170 , core_csr_decoded_decoded_andMatrixInput_2_171 }; 
    wire[5:0] core_csr_decoded_decoded_hi_171 ={ core_csr_decoded_decoded_hi_hi_171 , core_csr_decoded_decoded_hi_lo_170 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_163 ={ core_csr_decoded_decoded_andMatrixInput_9_171 , core_csr_decoded_decoded_andMatrixInput_10_170 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_171 ={ core_csr_decoded_decoded_lo_lo_hi_163 , core_csr_decoded_decoded_andMatrixInput_11_163 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_171 ={ core_csr_decoded_decoded_andMatrixInput_6_171 , core_csr_decoded_decoded_andMatrixInput_7_171 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_172 ={ core_csr_decoded_decoded_lo_hi_hi_171 , core_csr_decoded_decoded_andMatrixInput_8_171 }; 
    wire[5:0] core_csr_decoded_decoded_lo_172 ={ core_csr_decoded_decoded_lo_hi_172 , core_csr_decoded_decoded_lo_lo_171 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_170 ={ core_csr_decoded_decoded_andMatrixInput_3_172 , core_csr_decoded_decoded_andMatrixInput_4_172 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_171 ={ core_csr_decoded_decoded_hi_lo_hi_170 , core_csr_decoded_decoded_andMatrixInput_5_172 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_171 ={ core_csr_decoded_decoded_andMatrixInput_0_172 , core_csr_decoded_decoded_andMatrixInput_1_172 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_172 ={ core_csr_decoded_decoded_hi_hi_hi_171 , core_csr_decoded_decoded_andMatrixInput_2_172 }; 
    wire[5:0] core_csr_decoded_decoded_hi_172 ={ core_csr_decoded_decoded_hi_hi_172 , core_csr_decoded_decoded_hi_lo_171 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_164 ={ core_csr_decoded_decoded_andMatrixInput_9_172 , core_csr_decoded_decoded_andMatrixInput_10_171 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_172 ={ core_csr_decoded_decoded_lo_lo_hi_164 , core_csr_decoded_decoded_andMatrixInput_11_164 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_172 ={ core_csr_decoded_decoded_andMatrixInput_6_172 , core_csr_decoded_decoded_andMatrixInput_7_172 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_173 ={ core_csr_decoded_decoded_lo_hi_hi_172 , core_csr_decoded_decoded_andMatrixInput_8_172 }; 
    wire[5:0] core_csr_decoded_decoded_lo_173 ={ core_csr_decoded_decoded_lo_hi_173 , core_csr_decoded_decoded_lo_lo_172 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_171 ={ core_csr_decoded_decoded_andMatrixInput_3_173 , core_csr_decoded_decoded_andMatrixInput_4_173 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_172 ={ core_csr_decoded_decoded_hi_lo_hi_171 , core_csr_decoded_decoded_andMatrixInput_5_173 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_172 ={ core_csr_decoded_decoded_andMatrixInput_0_173 , core_csr_decoded_decoded_andMatrixInput_1_173 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_173 ={ core_csr_decoded_decoded_hi_hi_hi_172 , core_csr_decoded_decoded_andMatrixInput_2_173 }; 
    wire[5:0] core_csr_decoded_decoded_hi_173 ={ core_csr_decoded_decoded_hi_hi_173 , core_csr_decoded_decoded_hi_lo_172 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_165 ={ core_csr_decoded_decoded_andMatrixInput_9_173 , core_csr_decoded_decoded_andMatrixInput_10_172 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_173 ={ core_csr_decoded_decoded_lo_lo_hi_165 , core_csr_decoded_decoded_andMatrixInput_11_165 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_173 ={ core_csr_decoded_decoded_andMatrixInput_6_173 , core_csr_decoded_decoded_andMatrixInput_7_173 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_174 ={ core_csr_decoded_decoded_lo_hi_hi_173 , core_csr_decoded_decoded_andMatrixInput_8_173 }; 
    wire[5:0] core_csr_decoded_decoded_lo_174 ={ core_csr_decoded_decoded_lo_hi_174 , core_csr_decoded_decoded_lo_lo_173 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_172 ={ core_csr_decoded_decoded_andMatrixInput_3_174 , core_csr_decoded_decoded_andMatrixInput_4_174 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_173 ={ core_csr_decoded_decoded_hi_lo_hi_172 , core_csr_decoded_decoded_andMatrixInput_5_174 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_173 ={ core_csr_decoded_decoded_andMatrixInput_0_174 , core_csr_decoded_decoded_andMatrixInput_1_174 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_174 ={ core_csr_decoded_decoded_hi_hi_hi_173 , core_csr_decoded_decoded_andMatrixInput_2_174 }; 
    wire[5:0] core_csr_decoded_decoded_hi_174 ={ core_csr_decoded_decoded_hi_hi_174 , core_csr_decoded_decoded_hi_lo_173 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_166 ={ core_csr_decoded_decoded_andMatrixInput_9_174 , core_csr_decoded_decoded_andMatrixInput_10_173 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_174 ={ core_csr_decoded_decoded_lo_lo_hi_166 , core_csr_decoded_decoded_andMatrixInput_11_166 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_174 ={ core_csr_decoded_decoded_andMatrixInput_6_174 , core_csr_decoded_decoded_andMatrixInput_7_174 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_175 ={ core_csr_decoded_decoded_lo_hi_hi_174 , core_csr_decoded_decoded_andMatrixInput_8_174 }; 
    wire[5:0] core_csr_decoded_decoded_lo_175 ={ core_csr_decoded_decoded_lo_hi_175 , core_csr_decoded_decoded_lo_lo_174 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_173 ={ core_csr_decoded_decoded_andMatrixInput_3_175 , core_csr_decoded_decoded_andMatrixInput_4_175 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_174 ={ core_csr_decoded_decoded_hi_lo_hi_173 , core_csr_decoded_decoded_andMatrixInput_5_175 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_174 ={ core_csr_decoded_decoded_andMatrixInput_0_175 , core_csr_decoded_decoded_andMatrixInput_1_175 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_175 ={ core_csr_decoded_decoded_hi_hi_hi_174 , core_csr_decoded_decoded_andMatrixInput_2_175 }; 
    wire[5:0] core_csr_decoded_decoded_hi_175 ={ core_csr_decoded_decoded_hi_hi_175 , core_csr_decoded_decoded_hi_lo_174 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_167 ={ core_csr_decoded_decoded_andMatrixInput_9_175 , core_csr_decoded_decoded_andMatrixInput_10_174 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_175 ={ core_csr_decoded_decoded_lo_lo_hi_167 , core_csr_decoded_decoded_andMatrixInput_11_167 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_175 ={ core_csr_decoded_decoded_andMatrixInput_6_175 , core_csr_decoded_decoded_andMatrixInput_7_175 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_176 ={ core_csr_decoded_decoded_lo_hi_hi_175 , core_csr_decoded_decoded_andMatrixInput_8_175 }; 
    wire[5:0] core_csr_decoded_decoded_lo_176 ={ core_csr_decoded_decoded_lo_hi_176 , core_csr_decoded_decoded_lo_lo_175 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_174 ={ core_csr_decoded_decoded_andMatrixInput_3_176 , core_csr_decoded_decoded_andMatrixInput_4_176 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_175 ={ core_csr_decoded_decoded_hi_lo_hi_174 , core_csr_decoded_decoded_andMatrixInput_5_176 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_175 ={ core_csr_decoded_decoded_andMatrixInput_0_176 , core_csr_decoded_decoded_andMatrixInput_1_176 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_176 ={ core_csr_decoded_decoded_hi_hi_hi_175 , core_csr_decoded_decoded_andMatrixInput_2_176 }; 
    wire[5:0] core_csr_decoded_decoded_hi_176 ={ core_csr_decoded_decoded_hi_hi_176 , core_csr_decoded_decoded_hi_lo_175 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_168 ={ core_csr_decoded_decoded_andMatrixInput_9_176 , core_csr_decoded_decoded_andMatrixInput_10_175 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_176 ={ core_csr_decoded_decoded_lo_lo_hi_168 , core_csr_decoded_decoded_andMatrixInput_11_168 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_176 ={ core_csr_decoded_decoded_andMatrixInput_6_176 , core_csr_decoded_decoded_andMatrixInput_7_176 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_177 ={ core_csr_decoded_decoded_lo_hi_hi_176 , core_csr_decoded_decoded_andMatrixInput_8_176 }; 
    wire[5:0] core_csr_decoded_decoded_lo_177 ={ core_csr_decoded_decoded_lo_hi_177 , core_csr_decoded_decoded_lo_lo_176 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_175 ={ core_csr_decoded_decoded_andMatrixInput_3_177 , core_csr_decoded_decoded_andMatrixInput_4_177 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_176 ={ core_csr_decoded_decoded_hi_lo_hi_175 , core_csr_decoded_decoded_andMatrixInput_5_177 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_176 ={ core_csr_decoded_decoded_andMatrixInput_0_177 , core_csr_decoded_decoded_andMatrixInput_1_177 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_177 ={ core_csr_decoded_decoded_hi_hi_hi_176 , core_csr_decoded_decoded_andMatrixInput_2_177 }; 
    wire[5:0] core_csr_decoded_decoded_hi_177 ={ core_csr_decoded_decoded_hi_hi_177 , core_csr_decoded_decoded_hi_lo_176 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_169 ={ core_csr_decoded_decoded_andMatrixInput_9_177 , core_csr_decoded_decoded_andMatrixInput_10_176 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_177 ={ core_csr_decoded_decoded_lo_lo_hi_169 , core_csr_decoded_decoded_andMatrixInput_11_169 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_177 ={ core_csr_decoded_decoded_andMatrixInput_6_177 , core_csr_decoded_decoded_andMatrixInput_7_177 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_178 ={ core_csr_decoded_decoded_lo_hi_hi_177 , core_csr_decoded_decoded_andMatrixInput_8_177 }; 
    wire[5:0] core_csr_decoded_decoded_lo_178 ={ core_csr_decoded_decoded_lo_hi_178 , core_csr_decoded_decoded_lo_lo_177 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_176 ={ core_csr_decoded_decoded_andMatrixInput_3_178 , core_csr_decoded_decoded_andMatrixInput_4_178 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_177 ={ core_csr_decoded_decoded_hi_lo_hi_176 , core_csr_decoded_decoded_andMatrixInput_5_178 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_177 ={ core_csr_decoded_decoded_andMatrixInput_0_178 , core_csr_decoded_decoded_andMatrixInput_1_178 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_178 ={ core_csr_decoded_decoded_hi_hi_hi_177 , core_csr_decoded_decoded_andMatrixInput_2_178 }; 
    wire[5:0] core_csr_decoded_decoded_hi_178 ={ core_csr_decoded_decoded_hi_hi_178 , core_csr_decoded_decoded_hi_lo_177 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_170 ={ core_csr_decoded_decoded_andMatrixInput_9_178 , core_csr_decoded_decoded_andMatrixInput_10_177 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_178 ={ core_csr_decoded_decoded_lo_lo_hi_170 , core_csr_decoded_decoded_andMatrixInput_11_170 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_178 ={ core_csr_decoded_decoded_andMatrixInput_6_178 , core_csr_decoded_decoded_andMatrixInput_7_178 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_179 ={ core_csr_decoded_decoded_lo_hi_hi_178 , core_csr_decoded_decoded_andMatrixInput_8_178 }; 
    wire[5:0] core_csr_decoded_decoded_lo_179 ={ core_csr_decoded_decoded_lo_hi_179 , core_csr_decoded_decoded_lo_lo_178 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_177 ={ core_csr_decoded_decoded_andMatrixInput_3_179 , core_csr_decoded_decoded_andMatrixInput_4_179 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_178 ={ core_csr_decoded_decoded_hi_lo_hi_177 , core_csr_decoded_decoded_andMatrixInput_5_179 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_178 ={ core_csr_decoded_decoded_andMatrixInput_0_179 , core_csr_decoded_decoded_andMatrixInput_1_179 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_179 ={ core_csr_decoded_decoded_hi_hi_hi_178 , core_csr_decoded_decoded_andMatrixInput_2_179 }; 
    wire[5:0] core_csr_decoded_decoded_hi_179 ={ core_csr_decoded_decoded_hi_hi_179 , core_csr_decoded_decoded_hi_lo_178 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_171 ={ core_csr_decoded_decoded_andMatrixInput_9_179 , core_csr_decoded_decoded_andMatrixInput_10_178 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_179 ={ core_csr_decoded_decoded_lo_lo_hi_171 , core_csr_decoded_decoded_andMatrixInput_11_171 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_179 ={ core_csr_decoded_decoded_andMatrixInput_6_179 , core_csr_decoded_decoded_andMatrixInput_7_179 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_180 ={ core_csr_decoded_decoded_lo_hi_hi_179 , core_csr_decoded_decoded_andMatrixInput_8_179 }; 
    wire[5:0] core_csr_decoded_decoded_lo_180 ={ core_csr_decoded_decoded_lo_hi_180 , core_csr_decoded_decoded_lo_lo_179 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_178 ={ core_csr_decoded_decoded_andMatrixInput_3_180 , core_csr_decoded_decoded_andMatrixInput_4_180 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_179 ={ core_csr_decoded_decoded_hi_lo_hi_178 , core_csr_decoded_decoded_andMatrixInput_5_180 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_179 ={ core_csr_decoded_decoded_andMatrixInput_0_180 , core_csr_decoded_decoded_andMatrixInput_1_180 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_180 ={ core_csr_decoded_decoded_hi_hi_hi_179 , core_csr_decoded_decoded_andMatrixInput_2_180 }; 
    wire[5:0] core_csr_decoded_decoded_hi_180 ={ core_csr_decoded_decoded_hi_hi_180 , core_csr_decoded_decoded_hi_lo_179 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_172 ={ core_csr_decoded_decoded_andMatrixInput_9_180 , core_csr_decoded_decoded_andMatrixInput_10_179 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_180 ={ core_csr_decoded_decoded_lo_lo_hi_172 , core_csr_decoded_decoded_andMatrixInput_11_172 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_180 ={ core_csr_decoded_decoded_andMatrixInput_6_180 , core_csr_decoded_decoded_andMatrixInput_7_180 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_181 ={ core_csr_decoded_decoded_lo_hi_hi_180 , core_csr_decoded_decoded_andMatrixInput_8_180 }; 
    wire[5:0] core_csr_decoded_decoded_lo_181 ={ core_csr_decoded_decoded_lo_hi_181 , core_csr_decoded_decoded_lo_lo_180 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_179 ={ core_csr_decoded_decoded_andMatrixInput_3_181 , core_csr_decoded_decoded_andMatrixInput_4_181 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_180 ={ core_csr_decoded_decoded_hi_lo_hi_179 , core_csr_decoded_decoded_andMatrixInput_5_181 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_180 ={ core_csr_decoded_decoded_andMatrixInput_0_181 , core_csr_decoded_decoded_andMatrixInput_1_181 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_181 ={ core_csr_decoded_decoded_hi_hi_hi_180 , core_csr_decoded_decoded_andMatrixInput_2_181 }; 
    wire[5:0] core_csr_decoded_decoded_hi_181 ={ core_csr_decoded_decoded_hi_hi_181 , core_csr_decoded_decoded_hi_lo_180 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_173 ={ core_csr_decoded_decoded_andMatrixInput_9_181 , core_csr_decoded_decoded_andMatrixInput_10_180 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_181 ={ core_csr_decoded_decoded_lo_lo_hi_173 , core_csr_decoded_decoded_andMatrixInput_11_173 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_181 ={ core_csr_decoded_decoded_andMatrixInput_6_181 , core_csr_decoded_decoded_andMatrixInput_7_181 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_182 ={ core_csr_decoded_decoded_lo_hi_hi_181 , core_csr_decoded_decoded_andMatrixInput_8_181 }; 
    wire[5:0] core_csr_decoded_decoded_lo_182 ={ core_csr_decoded_decoded_lo_hi_182 , core_csr_decoded_decoded_lo_lo_181 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_180 ={ core_csr_decoded_decoded_andMatrixInput_3_182 , core_csr_decoded_decoded_andMatrixInput_4_182 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_181 ={ core_csr_decoded_decoded_hi_lo_hi_180 , core_csr_decoded_decoded_andMatrixInput_5_182 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_181 ={ core_csr_decoded_decoded_andMatrixInput_0_182 , core_csr_decoded_decoded_andMatrixInput_1_182 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_182 ={ core_csr_decoded_decoded_hi_hi_hi_181 , core_csr_decoded_decoded_andMatrixInput_2_182 }; 
    wire[5:0] core_csr_decoded_decoded_hi_182 ={ core_csr_decoded_decoded_hi_hi_182 , core_csr_decoded_decoded_hi_lo_181 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_174 ={ core_csr_decoded_decoded_andMatrixInput_9_182 , core_csr_decoded_decoded_andMatrixInput_10_181 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_182 ={ core_csr_decoded_decoded_lo_lo_hi_174 , core_csr_decoded_decoded_andMatrixInput_11_174 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_182 ={ core_csr_decoded_decoded_andMatrixInput_6_182 , core_csr_decoded_decoded_andMatrixInput_7_182 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_183 ={ core_csr_decoded_decoded_lo_hi_hi_182 , core_csr_decoded_decoded_andMatrixInput_8_182 }; 
    wire[5:0] core_csr_decoded_decoded_lo_183 ={ core_csr_decoded_decoded_lo_hi_183 , core_csr_decoded_decoded_lo_lo_182 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_181 ={ core_csr_decoded_decoded_andMatrixInput_3_183 , core_csr_decoded_decoded_andMatrixInput_4_183 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_182 ={ core_csr_decoded_decoded_hi_lo_hi_181 , core_csr_decoded_decoded_andMatrixInput_5_183 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_182 ={ core_csr_decoded_decoded_andMatrixInput_0_183 , core_csr_decoded_decoded_andMatrixInput_1_183 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_183 ={ core_csr_decoded_decoded_hi_hi_hi_182 , core_csr_decoded_decoded_andMatrixInput_2_183 }; 
    wire[5:0] core_csr_decoded_decoded_hi_183 ={ core_csr_decoded_decoded_hi_hi_183 , core_csr_decoded_decoded_hi_lo_182 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_175 ={ core_csr_decoded_decoded_andMatrixInput_9_183 , core_csr_decoded_decoded_andMatrixInput_10_182 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_183 ={ core_csr_decoded_decoded_lo_lo_hi_175 , core_csr_decoded_decoded_andMatrixInput_11_175 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_183 ={ core_csr_decoded_decoded_andMatrixInput_6_183 , core_csr_decoded_decoded_andMatrixInput_7_183 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_184 ={ core_csr_decoded_decoded_lo_hi_hi_183 , core_csr_decoded_decoded_andMatrixInput_8_183 }; 
    wire[5:0] core_csr_decoded_decoded_lo_184 ={ core_csr_decoded_decoded_lo_hi_184 , core_csr_decoded_decoded_lo_lo_183 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_182 ={ core_csr_decoded_decoded_andMatrixInput_3_184 , core_csr_decoded_decoded_andMatrixInput_4_184 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_183 ={ core_csr_decoded_decoded_hi_lo_hi_182 , core_csr_decoded_decoded_andMatrixInput_5_184 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_183 ={ core_csr_decoded_decoded_andMatrixInput_0_184 , core_csr_decoded_decoded_andMatrixInput_1_184 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_184 ={ core_csr_decoded_decoded_hi_hi_hi_183 , core_csr_decoded_decoded_andMatrixInput_2_184 }; 
    wire[5:0] core_csr_decoded_decoded_hi_184 ={ core_csr_decoded_decoded_hi_hi_184 , core_csr_decoded_decoded_hi_lo_183 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_176 ={ core_csr_decoded_decoded_andMatrixInput_9_184 , core_csr_decoded_decoded_andMatrixInput_10_183 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_184 ={ core_csr_decoded_decoded_lo_lo_hi_176 , core_csr_decoded_decoded_andMatrixInput_11_176 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_184 ={ core_csr_decoded_decoded_andMatrixInput_6_184 , core_csr_decoded_decoded_andMatrixInput_7_184 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_185 ={ core_csr_decoded_decoded_lo_hi_hi_184 , core_csr_decoded_decoded_andMatrixInput_8_184 }; 
    wire[5:0] core_csr_decoded_decoded_lo_185 ={ core_csr_decoded_decoded_lo_hi_185 , core_csr_decoded_decoded_lo_lo_184 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_183 ={ core_csr_decoded_decoded_andMatrixInput_3_185 , core_csr_decoded_decoded_andMatrixInput_4_185 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_184 ={ core_csr_decoded_decoded_hi_lo_hi_183 , core_csr_decoded_decoded_andMatrixInput_5_185 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_184 ={ core_csr_decoded_decoded_andMatrixInput_0_185 , core_csr_decoded_decoded_andMatrixInput_1_185 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_185 ={ core_csr_decoded_decoded_hi_hi_hi_184 , core_csr_decoded_decoded_andMatrixInput_2_185 }; 
    wire[5:0] core_csr_decoded_decoded_hi_185 ={ core_csr_decoded_decoded_hi_hi_185 , core_csr_decoded_decoded_hi_lo_184 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_177 ={ core_csr_decoded_decoded_andMatrixInput_9_185 , core_csr_decoded_decoded_andMatrixInput_10_184 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_185 ={ core_csr_decoded_decoded_lo_lo_hi_177 , core_csr_decoded_decoded_andMatrixInput_11_177 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_185 ={ core_csr_decoded_decoded_andMatrixInput_6_185 , core_csr_decoded_decoded_andMatrixInput_7_185 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_186 ={ core_csr_decoded_decoded_lo_hi_hi_185 , core_csr_decoded_decoded_andMatrixInput_8_185 }; 
    wire[5:0] core_csr_decoded_decoded_lo_186 ={ core_csr_decoded_decoded_lo_hi_186 , core_csr_decoded_decoded_lo_lo_185 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_184 ={ core_csr_decoded_decoded_andMatrixInput_3_186 , core_csr_decoded_decoded_andMatrixInput_4_186 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_185 ={ core_csr_decoded_decoded_hi_lo_hi_184 , core_csr_decoded_decoded_andMatrixInput_5_186 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_185 ={ core_csr_decoded_decoded_andMatrixInput_0_186 , core_csr_decoded_decoded_andMatrixInput_1_186 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_186 ={ core_csr_decoded_decoded_hi_hi_hi_185 , core_csr_decoded_decoded_andMatrixInput_2_186 }; 
    wire[5:0] core_csr_decoded_decoded_hi_186 ={ core_csr_decoded_decoded_hi_hi_186 , core_csr_decoded_decoded_hi_lo_185 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_178 ={ core_csr_decoded_decoded_andMatrixInput_9_186 , core_csr_decoded_decoded_andMatrixInput_10_185 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_186 ={ core_csr_decoded_decoded_lo_lo_hi_178 , core_csr_decoded_decoded_andMatrixInput_11_178 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_186 ={ core_csr_decoded_decoded_andMatrixInput_6_186 , core_csr_decoded_decoded_andMatrixInput_7_186 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_187 ={ core_csr_decoded_decoded_lo_hi_hi_186 , core_csr_decoded_decoded_andMatrixInput_8_186 }; 
    wire[5:0] core_csr_decoded_decoded_lo_187 ={ core_csr_decoded_decoded_lo_hi_187 , core_csr_decoded_decoded_lo_lo_186 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_185 ={ core_csr_decoded_decoded_andMatrixInput_3_187 , core_csr_decoded_decoded_andMatrixInput_4_187 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_186 ={ core_csr_decoded_decoded_hi_lo_hi_185 , core_csr_decoded_decoded_andMatrixInput_5_187 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_186 ={ core_csr_decoded_decoded_andMatrixInput_0_187 , core_csr_decoded_decoded_andMatrixInput_1_187 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_187 ={ core_csr_decoded_decoded_hi_hi_hi_186 , core_csr_decoded_decoded_andMatrixInput_2_187 }; 
    wire[5:0] core_csr_decoded_decoded_hi_187 ={ core_csr_decoded_decoded_hi_hi_187 , core_csr_decoded_decoded_hi_lo_186 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_179 ={ core_csr_decoded_decoded_andMatrixInput_9_187 , core_csr_decoded_decoded_andMatrixInput_10_186 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_187 ={ core_csr_decoded_decoded_lo_lo_hi_179 , core_csr_decoded_decoded_andMatrixInput_11_179 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_187 ={ core_csr_decoded_decoded_andMatrixInput_6_187 , core_csr_decoded_decoded_andMatrixInput_7_187 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_188 ={ core_csr_decoded_decoded_lo_hi_hi_187 , core_csr_decoded_decoded_andMatrixInput_8_187 }; 
    wire[5:0] core_csr_decoded_decoded_lo_188 ={ core_csr_decoded_decoded_lo_hi_188 , core_csr_decoded_decoded_lo_lo_187 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_186 ={ core_csr_decoded_decoded_andMatrixInput_3_188 , core_csr_decoded_decoded_andMatrixInput_4_188 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_187 ={ core_csr_decoded_decoded_hi_lo_hi_186 , core_csr_decoded_decoded_andMatrixInput_5_188 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_187 ={ core_csr_decoded_decoded_andMatrixInput_0_188 , core_csr_decoded_decoded_andMatrixInput_1_188 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_188 ={ core_csr_decoded_decoded_hi_hi_hi_187 , core_csr_decoded_decoded_andMatrixInput_2_188 }; 
    wire[5:0] core_csr_decoded_decoded_hi_188 ={ core_csr_decoded_decoded_hi_hi_188 , core_csr_decoded_decoded_hi_lo_187 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_180 ={ core_csr_decoded_decoded_andMatrixInput_9_188 , core_csr_decoded_decoded_andMatrixInput_10_187 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_188 ={ core_csr_decoded_decoded_lo_lo_hi_180 , core_csr_decoded_decoded_andMatrixInput_11_180 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_188 ={ core_csr_decoded_decoded_andMatrixInput_6_188 , core_csr_decoded_decoded_andMatrixInput_7_188 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_189 ={ core_csr_decoded_decoded_lo_hi_hi_188 , core_csr_decoded_decoded_andMatrixInput_8_188 }; 
    wire[5:0] core_csr_decoded_decoded_lo_189 ={ core_csr_decoded_decoded_lo_hi_189 , core_csr_decoded_decoded_lo_lo_188 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_187 ={ core_csr_decoded_decoded_andMatrixInput_3_189 , core_csr_decoded_decoded_andMatrixInput_4_189 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_188 ={ core_csr_decoded_decoded_hi_lo_hi_187 , core_csr_decoded_decoded_andMatrixInput_5_189 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_188 ={ core_csr_decoded_decoded_andMatrixInput_0_189 , core_csr_decoded_decoded_andMatrixInput_1_189 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_189 ={ core_csr_decoded_decoded_hi_hi_hi_188 , core_csr_decoded_decoded_andMatrixInput_2_189 }; 
    wire[5:0] core_csr_decoded_decoded_hi_189 ={ core_csr_decoded_decoded_hi_hi_189 , core_csr_decoded_decoded_hi_lo_188 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_181 ={ core_csr_decoded_decoded_andMatrixInput_9_189 , core_csr_decoded_decoded_andMatrixInput_10_188 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_189 ={ core_csr_decoded_decoded_lo_lo_hi_181 , core_csr_decoded_decoded_andMatrixInput_11_181 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_189 ={ core_csr_decoded_decoded_andMatrixInput_6_189 , core_csr_decoded_decoded_andMatrixInput_7_189 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_190 ={ core_csr_decoded_decoded_lo_hi_hi_189 , core_csr_decoded_decoded_andMatrixInput_8_189 }; 
    wire[5:0] core_csr_decoded_decoded_lo_190 ={ core_csr_decoded_decoded_lo_hi_190 , core_csr_decoded_decoded_lo_lo_189 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_188 ={ core_csr_decoded_decoded_andMatrixInput_3_190 , core_csr_decoded_decoded_andMatrixInput_4_190 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_189 ={ core_csr_decoded_decoded_hi_lo_hi_188 , core_csr_decoded_decoded_andMatrixInput_5_190 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_189 ={ core_csr_decoded_decoded_andMatrixInput_0_190 , core_csr_decoded_decoded_andMatrixInput_1_190 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_190 ={ core_csr_decoded_decoded_hi_hi_hi_189 , core_csr_decoded_decoded_andMatrixInput_2_190 }; 
    wire[5:0] core_csr_decoded_decoded_hi_190 ={ core_csr_decoded_decoded_hi_hi_190 , core_csr_decoded_decoded_hi_lo_189 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_190 ={ core_csr_decoded_decoded_andMatrixInput_9_190 , core_csr_decoded_decoded_andMatrixInput_10_189 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_190 ={ core_csr_decoded_decoded_andMatrixInput_6_190 , core_csr_decoded_decoded_andMatrixInput_7_190 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_191 ={ core_csr_decoded_decoded_lo_hi_hi_190 , core_csr_decoded_decoded_andMatrixInput_8_190 }; 
    wire[4:0] core_csr_decoded_decoded_lo_191 ={ core_csr_decoded_decoded_lo_hi_191 , core_csr_decoded_decoded_lo_lo_190 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_189 ={ core_csr_decoded_decoded_andMatrixInput_3_191 , core_csr_decoded_decoded_andMatrixInput_4_191 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_190 ={ core_csr_decoded_decoded_hi_lo_hi_189 , core_csr_decoded_decoded_andMatrixInput_5_191 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_190 ={ core_csr_decoded_decoded_andMatrixInput_0_191 , core_csr_decoded_decoded_andMatrixInput_1_191 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_191 ={ core_csr_decoded_decoded_hi_hi_hi_190 , core_csr_decoded_decoded_andMatrixInput_2_191 }; 
    wire[5:0] core_csr_decoded_decoded_hi_191 ={ core_csr_decoded_decoded_hi_hi_191 , core_csr_decoded_decoded_hi_lo_190 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_182 ={ core_csr_decoded_decoded_andMatrixInput_9_191 , core_csr_decoded_decoded_andMatrixInput_10_190 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_191 ={ core_csr_decoded_decoded_lo_lo_hi_182 , core_csr_decoded_decoded_andMatrixInput_11_182 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_191 ={ core_csr_decoded_decoded_andMatrixInput_6_191 , core_csr_decoded_decoded_andMatrixInput_7_191 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_192 ={ core_csr_decoded_decoded_lo_hi_hi_191 , core_csr_decoded_decoded_andMatrixInput_8_191 }; 
    wire[5:0] core_csr_decoded_decoded_lo_192 ={ core_csr_decoded_decoded_lo_hi_192 , core_csr_decoded_decoded_lo_lo_191 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_190 ={ core_csr_decoded_decoded_andMatrixInput_3_192 , core_csr_decoded_decoded_andMatrixInput_4_192 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_191 ={ core_csr_decoded_decoded_hi_lo_hi_190 , core_csr_decoded_decoded_andMatrixInput_5_192 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_191 ={ core_csr_decoded_decoded_andMatrixInput_0_192 , core_csr_decoded_decoded_andMatrixInput_1_192 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_192 ={ core_csr_decoded_decoded_hi_hi_hi_191 , core_csr_decoded_decoded_andMatrixInput_2_192 }; 
    wire[5:0] core_csr_decoded_decoded_hi_192 ={ core_csr_decoded_decoded_hi_hi_192 , core_csr_decoded_decoded_hi_lo_191 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_183 ={ core_csr_decoded_decoded_andMatrixInput_9_192 , core_csr_decoded_decoded_andMatrixInput_10_191 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_192 ={ core_csr_decoded_decoded_lo_lo_hi_183 , core_csr_decoded_decoded_andMatrixInput_11_183 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_192 ={ core_csr_decoded_decoded_andMatrixInput_6_192 , core_csr_decoded_decoded_andMatrixInput_7_192 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_193 ={ core_csr_decoded_decoded_lo_hi_hi_192 , core_csr_decoded_decoded_andMatrixInput_8_192 }; 
    wire[5:0] core_csr_decoded_decoded_lo_193 ={ core_csr_decoded_decoded_lo_hi_193 , core_csr_decoded_decoded_lo_lo_192 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_191 ={ core_csr_decoded_decoded_andMatrixInput_3_193 , core_csr_decoded_decoded_andMatrixInput_4_193 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_192 ={ core_csr_decoded_decoded_hi_lo_hi_191 , core_csr_decoded_decoded_andMatrixInput_5_193 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_192 ={ core_csr_decoded_decoded_andMatrixInput_0_193 , core_csr_decoded_decoded_andMatrixInput_1_193 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_193 ={ core_csr_decoded_decoded_hi_hi_hi_192 , core_csr_decoded_decoded_andMatrixInput_2_193 }; 
    wire[5:0] core_csr_decoded_decoded_hi_193 ={ core_csr_decoded_decoded_hi_hi_193 , core_csr_decoded_decoded_hi_lo_192 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_184 ={ core_csr_decoded_decoded_andMatrixInput_9_193 , core_csr_decoded_decoded_andMatrixInput_10_192 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_193 ={ core_csr_decoded_decoded_lo_lo_hi_184 , core_csr_decoded_decoded_andMatrixInput_11_184 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_193 ={ core_csr_decoded_decoded_andMatrixInput_6_193 , core_csr_decoded_decoded_andMatrixInput_7_193 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_194 ={ core_csr_decoded_decoded_lo_hi_hi_193 , core_csr_decoded_decoded_andMatrixInput_8_193 }; 
    wire[5:0] core_csr_decoded_decoded_lo_194 ={ core_csr_decoded_decoded_lo_hi_194 , core_csr_decoded_decoded_lo_lo_193 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_192 ={ core_csr_decoded_decoded_andMatrixInput_3_194 , core_csr_decoded_decoded_andMatrixInput_4_194 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_193 ={ core_csr_decoded_decoded_hi_lo_hi_192 , core_csr_decoded_decoded_andMatrixInput_5_194 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_193 ={ core_csr_decoded_decoded_andMatrixInput_0_194 , core_csr_decoded_decoded_andMatrixInput_1_194 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_194 ={ core_csr_decoded_decoded_hi_hi_hi_193 , core_csr_decoded_decoded_andMatrixInput_2_194 }; 
    wire[5:0] core_csr_decoded_decoded_hi_194 ={ core_csr_decoded_decoded_hi_hi_194 , core_csr_decoded_decoded_hi_lo_193 }; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_185 ={ core_csr_decoded_decoded_andMatrixInput_9_194 , core_csr_decoded_decoded_andMatrixInput_10_193 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_194 ={ core_csr_decoded_decoded_lo_lo_hi_185 , core_csr_decoded_decoded_andMatrixInput_11_185 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_194 ={ core_csr_decoded_decoded_andMatrixInput_6_194 , core_csr_decoded_decoded_andMatrixInput_7_194 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_195 ={ core_csr_decoded_decoded_lo_hi_hi_194 , core_csr_decoded_decoded_andMatrixInput_8_194 }; 
    wire[5:0] core_csr_decoded_decoded_lo_195 ={ core_csr_decoded_decoded_lo_hi_195 , core_csr_decoded_decoded_lo_lo_194 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_193 ={ core_csr_decoded_decoded_andMatrixInput_3_195 , core_csr_decoded_decoded_andMatrixInput_4_195 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_194 ={ core_csr_decoded_decoded_hi_lo_hi_193 , core_csr_decoded_decoded_andMatrixInput_5_195 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_194 ={ core_csr_decoded_decoded_andMatrixInput_0_195 , core_csr_decoded_decoded_andMatrixInput_1_195 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_195 ={ core_csr_decoded_decoded_hi_hi_hi_194 , core_csr_decoded_decoded_andMatrixInput_2_195 }; 
    wire[5:0] core_csr_decoded_decoded_hi_195 ={ core_csr_decoded_decoded_hi_hi_195 , core_csr_decoded_decoded_hi_lo_194 }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_191 , core_csr_decoded_decoded_lo_191 },&{ core_csr_decoded_decoded_hi_193 , core_csr_decoded_decoded_lo_193 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_195 , core_csr_decoded_decoded_lo_195 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_58 , core_csr_decoded_decoded_lo_58 },&{ core_csr_decoded_decoded_hi_66 , core_csr_decoded_decoded_lo_66 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_192 , core_csr_decoded_decoded_lo_192 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_55 , core_csr_decoded_decoded_lo_55 },&{ core_csr_decoded_decoded_hi_56 , core_csr_decoded_decoded_lo_56 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_57 , core_csr_decoded_decoded_lo_57 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_52 , core_csr_decoded_decoded_lo_52 },&{ core_csr_decoded_decoded_hi_53 , core_csr_decoded_decoded_lo_53 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_54 , core_csr_decoded_decoded_lo_54 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_49 , core_csr_decoded_decoded_lo_49 },&{ core_csr_decoded_decoded_hi_50 , core_csr_decoded_decoded_lo_50 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_51 , core_csr_decoded_decoded_lo_51 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_46 , core_csr_decoded_decoded_lo_46 },&{ core_csr_decoded_decoded_hi_47 , core_csr_decoded_decoded_lo_47 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_48 , core_csr_decoded_decoded_lo_48 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_43 , core_csr_decoded_decoded_lo_43 },&{ core_csr_decoded_decoded_hi_44 , core_csr_decoded_decoded_lo_44 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_45 , core_csr_decoded_decoded_lo_45 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_40 , core_csr_decoded_decoded_lo_40 },&{ core_csr_decoded_decoded_hi_41 , core_csr_decoded_decoded_lo_41 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_42 , core_csr_decoded_decoded_lo_42 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_160 , core_csr_decoded_decoded_lo_160 },&{ core_csr_decoded_decoded_hi_161 , core_csr_decoded_decoded_lo_161 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_39 , core_csr_decoded_decoded_lo_39 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_130 , core_csr_decoded_decoded_lo_130 },&{ core_csr_decoded_decoded_hi_98 , core_csr_decoded_decoded_lo_98 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_99 , core_csr_decoded_decoded_lo_99 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_128 , core_csr_decoded_decoded_lo_128 },&{ core_csr_decoded_decoded_hi_190 , core_csr_decoded_decoded_lo_190 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_129 , core_csr_decoded_decoded_lo_129 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_33 , core_csr_decoded_decoded_lo_33 },&{ core_csr_decoded_decoded_hi_97 , core_csr_decoded_decoded_lo_97 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_159 , core_csr_decoded_decoded_lo_159 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_158 , core_csr_decoded_decoded_lo_158 },&{ core_csr_decoded_decoded_hi_127 , core_csr_decoded_decoded_lo_127 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_189 , core_csr_decoded_decoded_lo_189 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_188 , core_csr_decoded_decoded_lo_188 },&{ core_csr_decoded_decoded_hi_32 , core_csr_decoded_decoded_lo_32 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_96 , core_csr_decoded_decoded_lo_96 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_95 , core_csr_decoded_decoded_lo_95 },&{ core_csr_decoded_decoded_hi_157 , core_csr_decoded_decoded_lo_157 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_126 , core_csr_decoded_decoded_lo_126 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi_lo ={&{ core_csr_decoded_decoded_hi_187 , core_csr_decoded_decoded_lo_187 },&{ core_csr_decoded_decoded_hi_31 , core_csr_decoded_decoded_lo_31 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_156 , core_csr_decoded_decoded_lo_156 },&{ core_csr_decoded_decoded_hi_125 , core_csr_decoded_decoded_lo_125 }}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_186 , core_csr_decoded_decoded_lo_186 },&{ core_csr_decoded_decoded_hi_30 , core_csr_decoded_decoded_lo_30 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_94 , core_csr_decoded_decoded_lo_94 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_93 , core_csr_decoded_decoded_lo_93 },&{ core_csr_decoded_decoded_hi_155 , core_csr_decoded_decoded_lo_155 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_124 , core_csr_decoded_decoded_lo_124 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_123 , core_csr_decoded_decoded_lo_123 },&{ core_csr_decoded_decoded_hi_185 , core_csr_decoded_decoded_lo_185 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_29 , core_csr_decoded_decoded_lo_29 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_28 , core_csr_decoded_decoded_lo_28 },&{ core_csr_decoded_decoded_hi_92 , core_csr_decoded_decoded_lo_92 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_154 , core_csr_decoded_decoded_lo_154 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_153 , core_csr_decoded_decoded_lo_153 },&{ core_csr_decoded_decoded_hi_122 , core_csr_decoded_decoded_lo_122 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_184 , core_csr_decoded_decoded_lo_184 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_183 , core_csr_decoded_decoded_lo_183 },&{ core_csr_decoded_decoded_hi_27 , core_csr_decoded_decoded_lo_27 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_91 , core_csr_decoded_decoded_lo_91 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_90 , core_csr_decoded_decoded_lo_90 },&{ core_csr_decoded_decoded_hi_152 , core_csr_decoded_decoded_lo_152 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_121 , core_csr_decoded_decoded_lo_121 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_120 , core_csr_decoded_decoded_lo_120 },&{ core_csr_decoded_decoded_hi_182 , core_csr_decoded_decoded_lo_182 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_26 , core_csr_decoded_decoded_lo_26 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_25 , core_csr_decoded_decoded_lo_25 },&{ core_csr_decoded_decoded_hi_89 , core_csr_decoded_decoded_lo_89 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_151 , core_csr_decoded_decoded_lo_151 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_150 , core_csr_decoded_decoded_lo_150 },&{ core_csr_decoded_decoded_hi_119 , core_csr_decoded_decoded_lo_119 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_181 , core_csr_decoded_decoded_lo_181 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_180 , core_csr_decoded_decoded_lo_180 },&{ core_csr_decoded_decoded_hi_24 , core_csr_decoded_decoded_lo_24 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_88 , core_csr_decoded_decoded_lo_88 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_87 , core_csr_decoded_decoded_lo_87 },&{ core_csr_decoded_decoded_hi_149 , core_csr_decoded_decoded_lo_149 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_118 , core_csr_decoded_decoded_lo_118 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_117 , core_csr_decoded_decoded_lo_117 },&{ core_csr_decoded_decoded_hi_179 , core_csr_decoded_decoded_lo_179 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_23 , core_csr_decoded_decoded_lo_23 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_22 , core_csr_decoded_decoded_lo_22 },&{ core_csr_decoded_decoded_hi_86 , core_csr_decoded_decoded_lo_86 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_148 , core_csr_decoded_decoded_lo_148 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_147 , core_csr_decoded_decoded_lo_147 },&{ core_csr_decoded_decoded_hi_116 , core_csr_decoded_decoded_lo_116 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_178 , core_csr_decoded_decoded_lo_178 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi_lo ={&{ core_csr_decoded_decoded_hi_21 , core_csr_decoded_decoded_lo_21 },&{ core_csr_decoded_decoded_hi_85 , core_csr_decoded_decoded_lo_85 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_115 , core_csr_decoded_decoded_lo_115 },&{ core_csr_decoded_decoded_hi_177 , core_csr_decoded_decoded_lo_177 }}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo }; 
    wire[97:0] core_csr_decoded_decoded_orMatrixOutputs_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_20 , core_csr_decoded_decoded_lo_20 },&{ core_csr_decoded_decoded_hi_84 , core_csr_decoded_decoded_lo_84 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_146 , core_csr_decoded_decoded_lo_146 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_145 , core_csr_decoded_decoded_lo_145 },&{ core_csr_decoded_decoded_hi_114 , core_csr_decoded_decoded_lo_114 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_176 , core_csr_decoded_decoded_lo_176 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_175 , core_csr_decoded_decoded_lo_175 },&{ core_csr_decoded_decoded_hi_19 , core_csr_decoded_decoded_lo_19 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_83 , core_csr_decoded_decoded_lo_83 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_82 , core_csr_decoded_decoded_lo_82 },&{ core_csr_decoded_decoded_hi_144 , core_csr_decoded_decoded_lo_144 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_113 , core_csr_decoded_decoded_lo_113 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_112 , core_csr_decoded_decoded_lo_112 },&{ core_csr_decoded_decoded_hi_174 , core_csr_decoded_decoded_lo_174 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_18 , core_csr_decoded_decoded_lo_18 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_17 , core_csr_decoded_decoded_lo_17 },&{ core_csr_decoded_decoded_hi_81 , core_csr_decoded_decoded_lo_81 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_143 , core_csr_decoded_decoded_lo_143 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_142 , core_csr_decoded_decoded_lo_142 },&{ core_csr_decoded_decoded_hi_111 , core_csr_decoded_decoded_lo_111 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_173 , core_csr_decoded_decoded_lo_173 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_172 , core_csr_decoded_decoded_lo_172 },&{ core_csr_decoded_decoded_hi_16 , core_csr_decoded_decoded_lo_16 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_80 , core_csr_decoded_decoded_lo_80 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_79 , core_csr_decoded_decoded_lo_79 },&{ core_csr_decoded_decoded_hi_141 , core_csr_decoded_decoded_lo_141 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_110 , core_csr_decoded_decoded_lo_110 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_109 , core_csr_decoded_decoded_lo_109 },&{ core_csr_decoded_decoded_hi_171 , core_csr_decoded_decoded_lo_171 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_15 , core_csr_decoded_decoded_lo_15 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_14 , core_csr_decoded_decoded_lo_14 },&{ core_csr_decoded_decoded_hi_78 , core_csr_decoded_decoded_lo_78 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_140 , core_csr_decoded_decoded_lo_140 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_139 , core_csr_decoded_decoded_lo_139 },&{ core_csr_decoded_decoded_hi_108 , core_csr_decoded_decoded_lo_108 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_170 , core_csr_decoded_decoded_lo_170 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_169 , core_csr_decoded_decoded_lo_169 },&{ core_csr_decoded_decoded_hi_13 , core_csr_decoded_decoded_lo_13 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_77 , core_csr_decoded_decoded_lo_77 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_76 , core_csr_decoded_decoded_lo_76 },&{ core_csr_decoded_decoded_hi_138 , core_csr_decoded_decoded_lo_138 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_107 , core_csr_decoded_decoded_lo_107 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_106 , core_csr_decoded_decoded_lo_106 },&{ core_csr_decoded_decoded_hi_168 , core_csr_decoded_decoded_lo_168 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_12 , core_csr_decoded_decoded_lo_12 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi_lo ={&{ core_csr_decoded_decoded_hi_75 , core_csr_decoded_decoded_lo_75 },&{ core_csr_decoded_decoded_hi_137 , core_csr_decoded_decoded_lo_137 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_167 , core_csr_decoded_decoded_lo_167 },&{ core_csr_decoded_decoded_hi_11 , core_csr_decoded_decoded_lo_11 }}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_74 , core_csr_decoded_decoded_lo_74 },&{ core_csr_decoded_decoded_hi_136 , core_csr_decoded_decoded_lo_136 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_105 , core_csr_decoded_decoded_lo_105 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_104 , core_csr_decoded_decoded_lo_104 },&{ core_csr_decoded_decoded_hi_166 , core_csr_decoded_decoded_lo_166 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_10 , core_csr_decoded_decoded_lo_10 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_9 , core_csr_decoded_decoded_lo_9 },&{ core_csr_decoded_decoded_hi_73 , core_csr_decoded_decoded_lo_73 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_135 , core_csr_decoded_decoded_lo_135 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_134 , core_csr_decoded_decoded_lo_134 },&{ core_csr_decoded_decoded_hi_103 , core_csr_decoded_decoded_lo_103 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_165 , core_csr_decoded_decoded_lo_165 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_164 , core_csr_decoded_decoded_lo_164 },&{ core_csr_decoded_decoded_hi_8 , core_csr_decoded_decoded_lo_8 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_72 , core_csr_decoded_decoded_lo_72 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_71 , core_csr_decoded_decoded_lo_71 },&{ core_csr_decoded_decoded_hi_133 , core_csr_decoded_decoded_lo_133 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_102 , core_csr_decoded_decoded_lo_102 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_101 , core_csr_decoded_decoded_lo_101 },&{ core_csr_decoded_decoded_hi_163 , core_csr_decoded_decoded_lo_163 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_7 , core_csr_decoded_decoded_lo_7 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_6 , core_csr_decoded_decoded_lo_6 },&{ core_csr_decoded_decoded_hi_70 , core_csr_decoded_decoded_lo_70 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_132 , core_csr_decoded_decoded_lo_132 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_131 , core_csr_decoded_decoded_lo_131 },&{ core_csr_decoded_decoded_hi_100 , core_csr_decoded_decoded_lo_100 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_162 , core_csr_decoded_decoded_lo_162 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_68 , core_csr_decoded_decoded_lo_68 },&{ core_csr_decoded_decoded_hi_5 , core_csr_decoded_decoded_lo_5 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_69 , core_csr_decoded_decoded_lo_69 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_65 , core_csr_decoded_decoded_lo_65 },&{ core_csr_decoded_decoded_hi_4 , core_csr_decoded_decoded_lo_4 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_67 , core_csr_decoded_decoded_lo_67 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_194 , core_csr_decoded_decoded_lo_194 },&{ core_csr_decoded_decoded_hi_63 , core_csr_decoded_decoded_lo_63 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_hi_hi ,&{ core_csr_decoded_decoded_hi_64 , core_csr_decoded_decoded_lo_64 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_lo_hi ={&{ core_csr_decoded_decoded_hi_35 , core_csr_decoded_decoded_lo_35 },&{ core_csr_decoded_decoded_hi_37 , core_csr_decoded_decoded_lo_37 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_lo_hi ,&{ core_csr_decoded_decoded_hi_36 , core_csr_decoded_decoded_lo_36 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_hi_hi ={&{ core_csr_decoded_decoded_hi_38 , core_csr_decoded_decoded_lo_38 },&{ core_csr_decoded_decoded_hi_2 , core_csr_decoded_decoded_lo_2 }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_hi_hi ,&{ core_csr_decoded_decoded_hi_34 , core_csr_decoded_decoded_lo_34 }}; 
    wire[5:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_lo_hi ={&{ core_csr_decoded_decoded_hi_1 , core_csr_decoded_decoded_lo_1 },&{ core_csr_decoded_decoded_hi , core_csr_decoded_decoded_lo }}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_lo_hi ,&{ core_csr_decoded_decoded_hi_3 , core_csr_decoded_decoded_lo_3 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi_lo ={&{ core_csr_decoded_decoded_hi_61 , core_csr_decoded_decoded_lo_61 },&{ core_csr_decoded_decoded_hi_62 , core_csr_decoded_decoded_lo_62 }}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi_hi ={&{ core_csr_decoded_decoded_hi_59 , core_csr_decoded_decoded_lo_59 },&{ core_csr_decoded_decoded_hi_60 , core_csr_decoded_decoded_lo_60 }}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo }; 
    wire[97:0] core_csr_decoded_decoded_orMatrixOutputs_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo }; 
    wire[195:0] core_csr_decoded_decoded_orMatrixOutputs ={ core_csr_decoded_decoded_orMatrixOutputs_hi , core_csr_decoded_decoded_orMatrixOutputs_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [2:1]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [0]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [5:4]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [3]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [8:7]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [6]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [11:10]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [9]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [14:13]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [12]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [17:16]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [15]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [20:19]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [18]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [23:22]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [21]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [26:25]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [24]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [29:28]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [27]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [32:31]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [30]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [35:34]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [33]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [38:37]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [36]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [41:40]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [39]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [44:43]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [42]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi_lo = core_csr_decoded_decoded_orMatrixOutputs [46:45]; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [48:47]; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [51:50]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [49]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [54:53]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [52]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [57:56]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [55]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [60:59]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [58]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [63:62]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [61]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [66:65]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [64]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [69:68]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [67]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [72:71]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [70]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [75:74]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [73]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [78:77]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [76]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [81:80]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [79]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [84:83]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [82]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [87:86]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [85]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [90:89]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [88]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [93:92]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [91]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi_lo = core_csr_decoded_decoded_orMatrixOutputs [95:94]; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [97:96]; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo }; 
    wire[97:0] core_csr_decoded_decoded_invMatrixOutputs_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [100:99]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [98]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [103:102]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [101]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [106:105]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [104]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [109:108]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [107]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [112:111]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [110]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [115:114]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [113]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [118:117]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [116]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [121:120]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [119]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [124:123]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [122]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [127:126]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [125]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [130:129]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [128]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [133:132]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [131]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [136:135]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [134]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [139:138]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [137]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [142:141]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [140]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi_lo = core_csr_decoded_decoded_orMatrixOutputs [144:143]; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [146:145]; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [149:148]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [147]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [152:151]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [150]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [155:154]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [153]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [158:157]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [156]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [161:160]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [159]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [164:163]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [162]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [167:166]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [165]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [170:169]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [168]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo }; 
    wire[23:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [173:172]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [171]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [176:175]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [174]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [179:178]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [177]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [182:181]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [180]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_lo }; 
    wire[11:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [185:184]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [183]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [188:187]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [186]}; 
    wire[5:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_lo_hi = core_csr_decoded_decoded_orMatrixOutputs [191:190]; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs [189]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi_lo = core_csr_decoded_decoded_orMatrixOutputs [193:192]; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi_hi = core_csr_decoded_decoded_orMatrixOutputs [195:194]; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi_lo }; 
    wire[6:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_lo }; 
    wire[12:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo }; 
    wire[24:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo }; 
    wire[48:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo }; 
    wire[97:0] core_csr_decoded_decoded_invMatrixOutputs_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo }; 
  assign  core_csr_decoded_decoded_invMatrixOutputs ={ core_csr_decoded_decoded_invMatrixOutputs_hi , core_csr_decoded_decoded_invMatrixOutputs_lo }; 
    wire[195:0] core_csr_decoded_decoded = core_csr_decoded_decoded_invMatrixOutputs ; 
  assign  core_csr_decoded_decoded_plaInput = core_csr_addr [11:0]; 
    wire core_csr_decoded_0 = core_csr_decoded_decoded [195]; 
    wire core_csr_decoded_1 = core_csr_decoded_decoded [194]; 
    wire core_csr_decoded_2 = core_csr_decoded_decoded [193]; 
    wire core_csr_decoded_3 = core_csr_decoded_decoded [192]; 
    wire core_csr_decoded_4 = core_csr_decoded_decoded [191]; 
    wire core_csr_decoded_5 = core_csr_decoded_decoded [190]; 
    wire core_csr_decoded_6 = core_csr_decoded_decoded [189]; 
    wire core_csr_decoded_7 = core_csr_decoded_decoded [188]; 
    wire core_csr_decoded_8 = core_csr_decoded_decoded [187]; 
    wire core_csr_decoded_9 = core_csr_decoded_decoded [186]; 
    wire core_csr_decoded_10 = core_csr_decoded_decoded [185]; 
    wire core_csr_decoded_11 = core_csr_decoded_decoded [184]; 
    wire core_csr_decoded_12 = core_csr_decoded_decoded [183]; 
    wire core_csr_decoded_13 = core_csr_decoded_decoded [182]; 
    wire core_csr_decoded_14 = core_csr_decoded_decoded [181]; 
    wire core_csr_decoded_15 = core_csr_decoded_decoded [180]; 
    wire core_csr_decoded_16 = core_csr_decoded_decoded [179]; 
    wire core_csr_decoded_17 = core_csr_decoded_decoded [178]; 
    wire core_csr_decoded_18 = core_csr_decoded_decoded [177]; 
    wire core_csr_decoded_19 = core_csr_decoded_decoded [176]; 
    wire core_csr_decoded_20 = core_csr_decoded_decoded [175]; 
    wire core_csr_decoded_21 = core_csr_decoded_decoded [174]; 
    wire core_csr_decoded_22 = core_csr_decoded_decoded [173]; 
    wire core_csr_decoded_23 = core_csr_decoded_decoded [172]; 
    wire core_csr_decoded_24 = core_csr_decoded_decoded [171]; 
    wire core_csr_decoded_25 = core_csr_decoded_decoded [170]; 
    wire core_csr_decoded_26 = core_csr_decoded_decoded [169]; 
    wire core_csr_decoded_27 = core_csr_decoded_decoded [168]; 
    wire core_csr_decoded_28 = core_csr_decoded_decoded [167]; 
    wire core_csr_decoded_29 = core_csr_decoded_decoded [166]; 
    wire core_csr_decoded_30 = core_csr_decoded_decoded [165]; 
    wire core_csr_decoded_31 = core_csr_decoded_decoded [164]; 
    wire core_csr_decoded_32 = core_csr_decoded_decoded [163]; 
    wire core_csr_decoded_33 = core_csr_decoded_decoded [162]; 
    wire core_csr_decoded_34 = core_csr_decoded_decoded [161]; 
    wire core_csr_decoded_35 = core_csr_decoded_decoded [160]; 
    wire core_csr_decoded_36 = core_csr_decoded_decoded [159]; 
    wire core_csr_decoded_37 = core_csr_decoded_decoded [158]; 
    wire core_csr_decoded_38 = core_csr_decoded_decoded [157]; 
    wire core_csr_decoded_39 = core_csr_decoded_decoded [156]; 
    wire core_csr_decoded_40 = core_csr_decoded_decoded [155]; 
    wire core_csr_decoded_41 = core_csr_decoded_decoded [154]; 
    wire core_csr_decoded_42 = core_csr_decoded_decoded [153]; 
    wire core_csr_decoded_43 = core_csr_decoded_decoded [152]; 
    wire core_csr_decoded_44 = core_csr_decoded_decoded [151]; 
    wire core_csr_decoded_45 = core_csr_decoded_decoded [150]; 
    wire core_csr_decoded_46 = core_csr_decoded_decoded [149]; 
    wire core_csr_decoded_47 = core_csr_decoded_decoded [148]; 
    wire core_csr_decoded_48 = core_csr_decoded_decoded [147]; 
    wire core_csr_decoded_49 = core_csr_decoded_decoded [146]; 
    wire core_csr_decoded_50 = core_csr_decoded_decoded [145]; 
    wire core_csr_decoded_51 = core_csr_decoded_decoded [144]; 
    wire core_csr_decoded_52 = core_csr_decoded_decoded [143]; 
    wire core_csr_decoded_53 = core_csr_decoded_decoded [142]; 
    wire core_csr_decoded_54 = core_csr_decoded_decoded [141]; 
    wire core_csr_decoded_55 = core_csr_decoded_decoded [140]; 
    wire core_csr_decoded_56 = core_csr_decoded_decoded [139]; 
    wire core_csr_decoded_57 = core_csr_decoded_decoded [138]; 
    wire core_csr_decoded_58 = core_csr_decoded_decoded [137]; 
    wire core_csr_decoded_59 = core_csr_decoded_decoded [136]; 
    wire core_csr_decoded_60 = core_csr_decoded_decoded [135]; 
    wire core_csr_decoded_61 = core_csr_decoded_decoded [134]; 
    wire core_csr_decoded_62 = core_csr_decoded_decoded [133]; 
    wire core_csr_decoded_63 = core_csr_decoded_decoded [132]; 
    wire core_csr_decoded_64 = core_csr_decoded_decoded [131]; 
    wire core_csr_decoded_65 = core_csr_decoded_decoded [130]; 
    wire core_csr_decoded_66 = core_csr_decoded_decoded [129]; 
    wire core_csr_decoded_67 = core_csr_decoded_decoded [128]; 
    wire core_csr_decoded_68 = core_csr_decoded_decoded [127]; 
    wire core_csr_decoded_69 = core_csr_decoded_decoded [126]; 
    wire core_csr_decoded_70 = core_csr_decoded_decoded [125]; 
    wire core_csr_decoded_71 = core_csr_decoded_decoded [124]; 
    wire core_csr_decoded_72 = core_csr_decoded_decoded [123]; 
    wire core_csr_decoded_73 = core_csr_decoded_decoded [122]; 
    wire core_csr_decoded_74 = core_csr_decoded_decoded [121]; 
    wire core_csr_decoded_75 = core_csr_decoded_decoded [120]; 
    wire core_csr_decoded_76 = core_csr_decoded_decoded [119]; 
    wire core_csr_decoded_77 = core_csr_decoded_decoded [118]; 
    wire core_csr_decoded_78 = core_csr_decoded_decoded [117]; 
    wire core_csr_decoded_79 = core_csr_decoded_decoded [116]; 
    wire core_csr_decoded_80 = core_csr_decoded_decoded [115]; 
    wire core_csr_decoded_81 = core_csr_decoded_decoded [114]; 
    wire core_csr_decoded_82 = core_csr_decoded_decoded [113]; 
    wire core_csr_decoded_83 = core_csr_decoded_decoded [112]; 
    wire core_csr_decoded_84 = core_csr_decoded_decoded [111]; 
    wire core_csr_decoded_85 = core_csr_decoded_decoded [110]; 
    wire core_csr_decoded_86 = core_csr_decoded_decoded [109]; 
    wire core_csr_decoded_87 = core_csr_decoded_decoded [108]; 
    wire core_csr_decoded_88 = core_csr_decoded_decoded [107]; 
    wire core_csr_decoded_89 = core_csr_decoded_decoded [106]; 
    wire core_csr_decoded_90 = core_csr_decoded_decoded [105]; 
    wire core_csr_decoded_91 = core_csr_decoded_decoded [104]; 
    wire core_csr_decoded_92 = core_csr_decoded_decoded [103]; 
    wire core_csr_decoded_93 = core_csr_decoded_decoded [102]; 
    wire core_csr_decoded_94 = core_csr_decoded_decoded [101]; 
    wire core_csr_decoded_95 = core_csr_decoded_decoded [100]; 
    wire core_csr_decoded_96 = core_csr_decoded_decoded [99]; 
    wire core_csr_decoded_97 = core_csr_decoded_decoded [98]; 
    wire core_csr_decoded_98 = core_csr_decoded_decoded [97]; 
    wire core_csr_decoded_99 = core_csr_decoded_decoded [96]; 
    wire core_csr_decoded_100 = core_csr_decoded_decoded [95]; 
    wire core_csr_decoded_101 = core_csr_decoded_decoded [94]; 
    wire core_csr_decoded_102 = core_csr_decoded_decoded [93]; 
    wire core_csr_decoded_103 = core_csr_decoded_decoded [92]; 
    wire core_csr_decoded_104 = core_csr_decoded_decoded [91]; 
    wire core_csr_decoded_105 = core_csr_decoded_decoded [90]; 
    wire core_csr_decoded_106 = core_csr_decoded_decoded [89]; 
    wire core_csr_decoded_107 = core_csr_decoded_decoded [88]; 
    wire core_csr_decoded_108 = core_csr_decoded_decoded [87]; 
    wire core_csr_decoded_109 = core_csr_decoded_decoded [86]; 
    wire core_csr_decoded_110 = core_csr_decoded_decoded [85]; 
    wire core_csr_decoded_111 = core_csr_decoded_decoded [84]; 
    wire core_csr_decoded_112 = core_csr_decoded_decoded [83]; 
    wire core_csr_decoded_113 = core_csr_decoded_decoded [82]; 
    wire core_csr_decoded_114 = core_csr_decoded_decoded [81]; 
    wire core_csr_decoded_115 = core_csr_decoded_decoded [80]; 
    wire core_csr_decoded_116 = core_csr_decoded_decoded [79]; 
    wire core_csr_decoded_117 = core_csr_decoded_decoded [78]; 
    wire core_csr_decoded_118 = core_csr_decoded_decoded [77]; 
    wire core_csr_decoded_119 = core_csr_decoded_decoded [76]; 
    wire core_csr_decoded_120 = core_csr_decoded_decoded [75]; 
    wire core_csr_decoded_121 = core_csr_decoded_decoded [74]; 
    wire core_csr_decoded_122 = core_csr_decoded_decoded [73]; 
    wire core_csr_decoded_123 = core_csr_decoded_decoded [72]; 
    wire core_csr_decoded_124 = core_csr_decoded_decoded [71]; 
    wire core_csr_decoded_125 = core_csr_decoded_decoded [70]; 
    wire core_csr_decoded_126 = core_csr_decoded_decoded [69]; 
    wire core_csr_decoded_127 = core_csr_decoded_decoded [68]; 
    wire core_csr_decoded_128 = core_csr_decoded_decoded [67]; 
    wire core_csr_decoded_129 = core_csr_decoded_decoded [66]; 
    wire core_csr_decoded_130 = core_csr_decoded_decoded [65]; 
    wire core_csr_decoded_131 = core_csr_decoded_decoded [64]; 
    wire core_csr_decoded_132 = core_csr_decoded_decoded [63]; 
    wire core_csr_decoded_133 = core_csr_decoded_decoded [62]; 
    wire core_csr_decoded_134 = core_csr_decoded_decoded [61]; 
    wire core_csr_decoded_135 = core_csr_decoded_decoded [60]; 
    wire core_csr_decoded_136 = core_csr_decoded_decoded [59]; 
    wire core_csr_decoded_137 = core_csr_decoded_decoded [58]; 
    wire core_csr_decoded_138 = core_csr_decoded_decoded [57]; 
    wire core_csr_decoded_139 = core_csr_decoded_decoded [56]; 
    wire core_csr_decoded_140 = core_csr_decoded_decoded [55]; 
    wire core_csr_decoded_141 = core_csr_decoded_decoded [54]; 
    wire core_csr_decoded_142 = core_csr_decoded_decoded [53]; 
    wire core_csr_decoded_143 = core_csr_decoded_decoded [52]; 
    wire core_csr_decoded_144 = core_csr_decoded_decoded [51]; 
    wire core_csr_decoded_145 = core_csr_decoded_decoded [50]; 
    wire core_csr_decoded_146 = core_csr_decoded_decoded [49]; 
    wire core_csr_decoded_147 = core_csr_decoded_decoded [48]; 
    wire core_csr_decoded_148 = core_csr_decoded_decoded [47]; 
    wire core_csr_decoded_149 = core_csr_decoded_decoded [46]; 
    wire core_csr_decoded_150 = core_csr_decoded_decoded [45]; 
    wire core_csr_decoded_151 = core_csr_decoded_decoded [44]; 
    wire core_csr_decoded_152 = core_csr_decoded_decoded [43]; 
    wire core_csr_decoded_153 = core_csr_decoded_decoded [42]; 
    wire core_csr_decoded_154 = core_csr_decoded_decoded [41]; 
    wire core_csr_decoded_155 = core_csr_decoded_decoded [40]; 
    wire core_csr_decoded_156 = core_csr_decoded_decoded [39]; 
    wire core_csr_decoded_157 = core_csr_decoded_decoded [38]; 
    wire core_csr_decoded_158 = core_csr_decoded_decoded [37]; 
    wire core_csr_decoded_159 = core_csr_decoded_decoded [36]; 
    wire core_csr_decoded_160 = core_csr_decoded_decoded [35]; 
    wire core_csr_decoded_161 = core_csr_decoded_decoded [34]; 
    wire core_csr_decoded_162 = core_csr_decoded_decoded [33]; 
    wire core_csr_decoded_163 = core_csr_decoded_decoded [32]; 
    wire core_csr_decoded_164 = core_csr_decoded_decoded [31]; 
    wire core_csr_decoded_165 = core_csr_decoded_decoded [30]; 
    wire core_csr_decoded_166 = core_csr_decoded_decoded [29]; 
    wire core_csr_decoded_167 = core_csr_decoded_decoded [28]; 
    wire core_csr_decoded_168 = core_csr_decoded_decoded [27]; 
    wire core_csr_decoded_169 = core_csr_decoded_decoded [26]; 
    wire core_csr_decoded_170 = core_csr_decoded_decoded [25]; 
    wire core_csr_decoded_171 = core_csr_decoded_decoded [24]; 
    wire core_csr_decoded_172 = core_csr_decoded_decoded [23]; 
    wire core_csr_decoded_173 = core_csr_decoded_decoded [22]; 
    wire core_csr_decoded_174 = core_csr_decoded_decoded [21]; 
    wire core_csr_decoded_175 = core_csr_decoded_decoded [20]; 
    wire core_csr_decoded_176 = core_csr_decoded_decoded [19]; 
    wire core_csr_decoded_177 = core_csr_decoded_decoded [18]; 
    wire core_csr_decoded_178 = core_csr_decoded_decoded [17]; 
    wire core_csr_decoded_179 = core_csr_decoded_decoded [16]; 
    wire core_csr_decoded_180 = core_csr_decoded_decoded [15]; 
    wire core_csr_decoded_181 = core_csr_decoded_decoded [14]; 
    wire core_csr_decoded_182 = core_csr_decoded_decoded [13]; 
    wire core_csr_decoded_183 = core_csr_decoded_decoded [12]; 
    wire core_csr_decoded_184 = core_csr_decoded_decoded [11]; 
    wire core_csr_decoded_185 = core_csr_decoded_decoded [10]; 
    wire core_csr_decoded_186 = core_csr_decoded_decoded [9]; 
    wire core_csr_decoded_187 = core_csr_decoded_decoded [8]; 
    wire core_csr_decoded_188 = core_csr_decoded_decoded [7]; 
    wire core_csr_decoded_189 = core_csr_decoded_decoded [6]; 
    wire core_csr_decoded_190 = core_csr_decoded_decoded [5]; 
    wire core_csr_decoded_191 = core_csr_decoded_decoded [4]; 
    wire core_csr_decoded_192 = core_csr_decoded_decoded [3]; 
    wire core_csr_decoded_193 = core_csr_decoded_decoded [2]; 
    wire core_csr_decoded_194 = core_csr_decoded_decoded [1]; 
    wire core_csr_decoded_195 = core_csr_decoded_decoded [0]; 
    wire[31:0] core_csr_wdata =(( core_csr_io_rw_cmd [1] ?  core_csr__io_rw_rdata_output :32'h0)| core_csr_io_rw_wdata )&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :32'h0); 
    wire core_csr_system_insn = core_csr_io_rw_cmd ==3'h4; 
    wire[31:0] core_csr_insn ={ core_csr_io_rw_addr ,20'h73}; 
    wire[31:0] core_csr_decoded_plaInput = core_csr_insn ; 
    wire[31:0] core_csr_decoded_invInputs =~ core_csr_decoded_plaInput ; 
    wire[8:0] core_csr_decoded_invMatrixOutputs ; 
    wire core_csr_decoded_andMatrixInput_0 = core_csr_decoded_invInputs [20]; 
    wire core_csr_decoded_andMatrixInput_1 = core_csr_decoded_invInputs [21]; 
    wire core_csr_decoded_andMatrixInput_1_1 = core_csr_decoded_invInputs [21]; 
    wire core_csr_decoded_andMatrixInput_2 = core_csr_decoded_invInputs [22]; 
    wire core_csr_decoded_andMatrixInput_2_1 = core_csr_decoded_invInputs [22]; 
    wire core_csr_decoded_andMatrixInput_0_3 = core_csr_decoded_invInputs [22]; 
    wire core_csr_decoded_andMatrixInput_3 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_3_1 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_1_3 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_1_4 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_4 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_4_1 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_2_3 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_2_4 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_5 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_5_1 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_3_3 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_3_4 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_6 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_6_1 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_4_2 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_4_3 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_7 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_7_1 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_5_2 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_5_3 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_8 = core_csr_decoded_invInputs [28]; 
    wire core_csr_decoded_andMatrixInput_8_1 = core_csr_decoded_invInputs [28]; 
    wire core_csr_decoded_andMatrixInput_9 = core_csr_decoded_invInputs [29]; 
    wire core_csr_decoded_andMatrixInput_9_1 = core_csr_decoded_invInputs [29]; 
    wire core_csr_decoded_andMatrixInput_1_2 = core_csr_decoded_invInputs [29]; 
    wire core_csr_decoded_andMatrixInput_10 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_10_1 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_2_2 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_8_2 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_8_3 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_11 = core_csr_decoded_invInputs [31]; 
    wire core_csr_decoded_andMatrixInput_11_1 = core_csr_decoded_invInputs [31]; 
    wire core_csr_decoded_andMatrixInput_3_2 = core_csr_decoded_invInputs [31]; 
    wire core_csr_decoded_andMatrixInput_9_2 = core_csr_decoded_invInputs [31]; 
    wire core_csr_decoded_andMatrixInput_9_3 = core_csr_decoded_invInputs [31]; 
    wire core_csr_decoded_andMatrixInput_1_5 = core_csr_decoded_invInputs [31]; 
    wire[1:0] core_csr_decoded_lo_lo_hi ={ core_csr_decoded_andMatrixInput_9 , core_csr_decoded_andMatrixInput_10 }; 
    wire[2:0] core_csr_decoded_lo_lo ={ core_csr_decoded_lo_lo_hi , core_csr_decoded_andMatrixInput_11 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi ={ core_csr_decoded_andMatrixInput_6 , core_csr_decoded_andMatrixInput_7 }; 
    wire[2:0] core_csr_decoded_lo_hi ={ core_csr_decoded_lo_hi_hi , core_csr_decoded_andMatrixInput_8 }; 
    wire[5:0] core_csr_decoded_lo ={ core_csr_decoded_lo_hi , core_csr_decoded_lo_lo }; 
    wire[1:0] core_csr_decoded_hi_lo_hi ={ core_csr_decoded_andMatrixInput_3 , core_csr_decoded_andMatrixInput_4 }; 
    wire[2:0] core_csr_decoded_hi_lo ={ core_csr_decoded_hi_lo_hi , core_csr_decoded_andMatrixInput_5 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi ={ core_csr_decoded_andMatrixInput_0 , core_csr_decoded_andMatrixInput_1 }; 
    wire[2:0] core_csr_decoded_hi_hi ={ core_csr_decoded_hi_hi_hi , core_csr_decoded_andMatrixInput_2 }; 
    wire[5:0] core_csr_decoded_hi ={ core_csr_decoded_hi_hi , core_csr_decoded_hi_lo }; 
    wire core_csr_decoded_andMatrixInput_0_1 = core_csr_decoded_plaInput [20]; 
    wire[1:0] core_csr_decoded_lo_lo_hi_1 ={ core_csr_decoded_andMatrixInput_9_1 , core_csr_decoded_andMatrixInput_10_1 }; 
    wire[2:0] core_csr_decoded_lo_lo_1 ={ core_csr_decoded_lo_lo_hi_1 , core_csr_decoded_andMatrixInput_11_1 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_1 ={ core_csr_decoded_andMatrixInput_6_1 , core_csr_decoded_andMatrixInput_7_1 }; 
    wire[2:0] core_csr_decoded_lo_hi_1 ={ core_csr_decoded_lo_hi_hi_1 , core_csr_decoded_andMatrixInput_8_1 }; 
    wire[5:0] core_csr_decoded_lo_1 ={ core_csr_decoded_lo_hi_1 , core_csr_decoded_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_hi_lo_hi_1 ={ core_csr_decoded_andMatrixInput_3_1 , core_csr_decoded_andMatrixInput_4_1 }; 
    wire[2:0] core_csr_decoded_hi_lo_1 ={ core_csr_decoded_hi_lo_hi_1 , core_csr_decoded_andMatrixInput_5_1 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_1 ={ core_csr_decoded_andMatrixInput_0_1 , core_csr_decoded_andMatrixInput_1_1 }; 
    wire[2:0] core_csr_decoded_hi_hi_1 ={ core_csr_decoded_hi_hi_hi_1 , core_csr_decoded_andMatrixInput_2_1 }; 
    wire[5:0] core_csr_decoded_hi_1 ={ core_csr_decoded_hi_hi_1 , core_csr_decoded_hi_lo_1 }; 
    wire core_csr_decoded_andMatrixInput_0_2 = core_csr_decoded_plaInput [28]; 
    wire core_csr_decoded_andMatrixInput_6_2 = core_csr_decoded_plaInput [28]; 
    wire core_csr_decoded_andMatrixInput_6_3 = core_csr_decoded_plaInput [28]; 
    wire[1:0] core_csr_decoded_lo_2 ={ core_csr_decoded_andMatrixInput_2_2 , core_csr_decoded_andMatrixInput_3_2 }; 
    wire[1:0] core_csr_decoded_hi_2 ={ core_csr_decoded_andMatrixInput_0_2 , core_csr_decoded_andMatrixInput_1_2 }; 
    wire core_csr_decoded_andMatrixInput_7_2 = core_csr_decoded_plaInput [29]; 
    wire core_csr_decoded_andMatrixInput_7_3 = core_csr_decoded_plaInput [29]; 
    wire[1:0] core_csr_decoded_lo_lo_2 ={ core_csr_decoded_andMatrixInput_8_2 , core_csr_decoded_andMatrixInput_9_2 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_2 ={ core_csr_decoded_andMatrixInput_5_2 , core_csr_decoded_andMatrixInput_6_2 }; 
    wire[2:0] core_csr_decoded_lo_hi_2 ={ core_csr_decoded_lo_hi_hi_2 , core_csr_decoded_andMatrixInput_7_2 }; 
    wire[4:0] core_csr_decoded_lo_3 ={ core_csr_decoded_lo_hi_2 , core_csr_decoded_lo_lo_2 }; 
    wire[1:0] core_csr_decoded_hi_lo_2 ={ core_csr_decoded_andMatrixInput_3_3 , core_csr_decoded_andMatrixInput_4_2 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_2 ={ core_csr_decoded_andMatrixInput_0_3 , core_csr_decoded_andMatrixInput_1_3 }; 
    wire[2:0] core_csr_decoded_hi_hi_2 ={ core_csr_decoded_hi_hi_hi_2 , core_csr_decoded_andMatrixInput_2_3 }; 
    wire[4:0] core_csr_decoded_hi_3 ={ core_csr_decoded_hi_hi_2 , core_csr_decoded_hi_lo_2 }; 
    wire core_csr_decoded_andMatrixInput_0_4 = core_csr_decoded_plaInput [22]; 
    wire[1:0] core_csr_decoded_lo_lo_3 ={ core_csr_decoded_andMatrixInput_8_3 , core_csr_decoded_andMatrixInput_9_3 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_3 ={ core_csr_decoded_andMatrixInput_5_3 , core_csr_decoded_andMatrixInput_6_3 }; 
    wire[2:0] core_csr_decoded_lo_hi_3 ={ core_csr_decoded_lo_hi_hi_3 , core_csr_decoded_andMatrixInput_7_3 }; 
    wire[4:0] core_csr_decoded_lo_4 ={ core_csr_decoded_lo_hi_3 , core_csr_decoded_lo_lo_3 }; 
    wire[1:0] core_csr_decoded_hi_lo_3 ={ core_csr_decoded_andMatrixInput_3_4 , core_csr_decoded_andMatrixInput_4_3 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_3 ={ core_csr_decoded_andMatrixInput_0_4 , core_csr_decoded_andMatrixInput_1_4 }; 
    wire[2:0] core_csr_decoded_hi_hi_3 ={ core_csr_decoded_hi_hi_hi_3 , core_csr_decoded_andMatrixInput_2_4 }; 
    wire[4:0] core_csr_decoded_hi_4 ={ core_csr_decoded_hi_hi_3 , core_csr_decoded_hi_lo_3 }; 
    wire core_csr_decoded_andMatrixInput_0_5 = core_csr_decoded_plaInput [30]; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_lo ={&{ core_csr_decoded_hi_4 , core_csr_decoded_lo_4 },&{ core_csr_decoded_hi_2 , core_csr_decoded_lo_2 }}; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_hi_hi ={&{ core_csr_decoded_hi , core_csr_decoded_lo },&{ core_csr_decoded_hi_1 , core_csr_decoded_lo_1 }}; 
    wire[2:0] core_csr_decoded_orMatrixOutputs_hi_hi ={ core_csr_decoded_orMatrixOutputs_hi_hi_hi ,|{&{ core_csr_decoded_hi_3 , core_csr_decoded_lo_3 },&{ core_csr_decoded_andMatrixInput_0_5 , core_csr_decoded_andMatrixInput_1_5 }}}; 
    wire[4:0] core_csr_decoded_orMatrixOutputs_hi ={ core_csr_decoded_orMatrixOutputs_hi_hi , core_csr_decoded_orMatrixOutputs_hi_lo }; 
    wire[8:0] core_csr_decoded_orMatrixOutputs ={ core_csr_decoded_orMatrixOutputs_hi ,4'h0}; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_lo = core_csr_decoded_orMatrixOutputs [1:0]; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_hi = core_csr_decoded_orMatrixOutputs [3:2]; 
    wire[3:0] core_csr_decoded_invMatrixOutputs_lo ={ core_csr_decoded_invMatrixOutputs_lo_hi , core_csr_decoded_invMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_lo = core_csr_decoded_orMatrixOutputs [5:4]; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_hi_hi = core_csr_decoded_orMatrixOutputs [8:7]; 
    wire[2:0] core_csr_decoded_invMatrixOutputs_hi_hi ={ core_csr_decoded_invMatrixOutputs_hi_hi_hi , core_csr_decoded_orMatrixOutputs [6]}; 
    wire[4:0] core_csr_decoded_invMatrixOutputs_hi ={ core_csr_decoded_invMatrixOutputs_hi_hi , core_csr_decoded_invMatrixOutputs_hi_lo }; 
  assign  core_csr_decoded_invMatrixOutputs ={ core_csr_decoded_invMatrixOutputs_hi , core_csr_decoded_invMatrixOutputs_lo }; 
    wire[8:0] core_csr_decoded = core_csr_decoded_invMatrixOutputs ; 
    wire core_csr_insn_call = core_csr_system_insn & core_csr_decoded [8]; 
    wire core_csr_insn_break = core_csr_system_insn & core_csr_decoded [7]; 
    wire core_csr_insn_ret = core_csr_system_insn & core_csr_decoded [6]; 
    wire core_csr_insn_cease = core_csr_system_insn & core_csr_decoded [5]; 
    wire core_csr_insn_wfi = core_csr_system_insn & core_csr_decoded [4]; 
    wire[11:0] core_csr_addr_1 = core_csr_io_decode_0_inst [31:20]; 
    wire[11:0] core_csr_io_decode_0_fp_csr_plaInput = core_csr_addr_1 ; 
    wire[11:0] core_csr_io_decode_0_read_illegal_plaInput = core_csr_addr_1 ; 
    wire[11:0] core_csr_io_decode_0_read_illegal_plaInput_1 = core_csr_addr_1 ; 
    wire[31:0] core_csr_decoded_invInputs_1 =~ core_csr_decoded_plaInput_1 ; 
    wire[8:0] core_csr_decoded_invMatrixOutputs_1 ; 
    wire core_csr_decoded_andMatrixInput_0_6 = core_csr_decoded_invInputs_1 [20]; 
    wire core_csr_decoded_andMatrixInput_1_6 = core_csr_decoded_invInputs_1 [21]; 
    wire core_csr_decoded_andMatrixInput_1_7 = core_csr_decoded_invInputs_1 [21]; 
    wire core_csr_decoded_andMatrixInput_2_5 = core_csr_decoded_invInputs_1 [22]; 
    wire core_csr_decoded_andMatrixInput_2_6 = core_csr_decoded_invInputs_1 [22]; 
    wire core_csr_decoded_andMatrixInput_0_9 = core_csr_decoded_invInputs_1 [22]; 
    wire core_csr_decoded_andMatrixInput_3_5 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_3_6 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_1_9 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_1_10 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_4_4 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_4_5 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_2_8 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_2_9 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_5_4 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_5_5 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_3_8 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_3_9 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_6_4 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_6_5 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_4_6 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_4_7 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_7_4 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_7_5 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_5_6 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_5_7 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_8_4 = core_csr_decoded_invInputs_1 [28]; 
    wire core_csr_decoded_andMatrixInput_8_5 = core_csr_decoded_invInputs_1 [28]; 
    wire core_csr_decoded_andMatrixInput_9_4 = core_csr_decoded_invInputs_1 [29]; 
    wire core_csr_decoded_andMatrixInput_9_5 = core_csr_decoded_invInputs_1 [29]; 
    wire core_csr_decoded_andMatrixInput_1_8 = core_csr_decoded_invInputs_1 [29]; 
    wire core_csr_decoded_andMatrixInput_10_2 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_10_3 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_2_7 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_8_6 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_8_7 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_11_2 = core_csr_decoded_invInputs_1 [31]; 
    wire core_csr_decoded_andMatrixInput_11_3 = core_csr_decoded_invInputs_1 [31]; 
    wire core_csr_decoded_andMatrixInput_3_7 = core_csr_decoded_invInputs_1 [31]; 
    wire core_csr_decoded_andMatrixInput_9_6 = core_csr_decoded_invInputs_1 [31]; 
    wire core_csr_decoded_andMatrixInput_9_7 = core_csr_decoded_invInputs_1 [31]; 
    wire core_csr_decoded_andMatrixInput_1_11 = core_csr_decoded_invInputs_1 [31]; 
    wire[1:0] core_csr_decoded_lo_lo_hi_2 ={ core_csr_decoded_andMatrixInput_9_4 , core_csr_decoded_andMatrixInput_10_2 }; 
    wire[2:0] core_csr_decoded_lo_lo_4 ={ core_csr_decoded_lo_lo_hi_2 , core_csr_decoded_andMatrixInput_11_2 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_4 ={ core_csr_decoded_andMatrixInput_6_4 , core_csr_decoded_andMatrixInput_7_4 }; 
    wire[2:0] core_csr_decoded_lo_hi_4 ={ core_csr_decoded_lo_hi_hi_4 , core_csr_decoded_andMatrixInput_8_4 }; 
    wire[5:0] core_csr_decoded_lo_5 ={ core_csr_decoded_lo_hi_4 , core_csr_decoded_lo_lo_4 }; 
    wire[1:0] core_csr_decoded_hi_lo_hi_2 ={ core_csr_decoded_andMatrixInput_3_5 , core_csr_decoded_andMatrixInput_4_4 }; 
    wire[2:0] core_csr_decoded_hi_lo_4 ={ core_csr_decoded_hi_lo_hi_2 , core_csr_decoded_andMatrixInput_5_4 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_4 ={ core_csr_decoded_andMatrixInput_0_6 , core_csr_decoded_andMatrixInput_1_6 }; 
    wire[2:0] core_csr_decoded_hi_hi_4 ={ core_csr_decoded_hi_hi_hi_4 , core_csr_decoded_andMatrixInput_2_5 }; 
    wire[5:0] core_csr_decoded_hi_5 ={ core_csr_decoded_hi_hi_4 , core_csr_decoded_hi_lo_4 }; 
    wire core_csr_decoded_andMatrixInput_0_7 = core_csr_decoded_plaInput_1 [20]; 
    wire[1:0] core_csr_decoded_lo_lo_hi_3 ={ core_csr_decoded_andMatrixInput_9_5 , core_csr_decoded_andMatrixInput_10_3 }; 
    wire[2:0] core_csr_decoded_lo_lo_5 ={ core_csr_decoded_lo_lo_hi_3 , core_csr_decoded_andMatrixInput_11_3 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_5 ={ core_csr_decoded_andMatrixInput_6_5 , core_csr_decoded_andMatrixInput_7_5 }; 
    wire[2:0] core_csr_decoded_lo_hi_5 ={ core_csr_decoded_lo_hi_hi_5 , core_csr_decoded_andMatrixInput_8_5 }; 
    wire[5:0] core_csr_decoded_lo_6 ={ core_csr_decoded_lo_hi_5 , core_csr_decoded_lo_lo_5 }; 
    wire[1:0] core_csr_decoded_hi_lo_hi_3 ={ core_csr_decoded_andMatrixInput_3_6 , core_csr_decoded_andMatrixInput_4_5 }; 
    wire[2:0] core_csr_decoded_hi_lo_5 ={ core_csr_decoded_hi_lo_hi_3 , core_csr_decoded_andMatrixInput_5_5 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_5 ={ core_csr_decoded_andMatrixInput_0_7 , core_csr_decoded_andMatrixInput_1_7 }; 
    wire[2:0] core_csr_decoded_hi_hi_5 ={ core_csr_decoded_hi_hi_hi_5 , core_csr_decoded_andMatrixInput_2_6 }; 
    wire[5:0] core_csr_decoded_hi_6 ={ core_csr_decoded_hi_hi_5 , core_csr_decoded_hi_lo_5 }; 
    wire core_csr_decoded_andMatrixInput_0_8 = core_csr_decoded_plaInput_1 [28]; 
    wire core_csr_decoded_andMatrixInput_6_6 = core_csr_decoded_plaInput_1 [28]; 
    wire core_csr_decoded_andMatrixInput_6_7 = core_csr_decoded_plaInput_1 [28]; 
    wire[1:0] core_csr_decoded_lo_7 ={ core_csr_decoded_andMatrixInput_2_7 , core_csr_decoded_andMatrixInput_3_7 }; 
    wire[1:0] core_csr_decoded_hi_7 ={ core_csr_decoded_andMatrixInput_0_8 , core_csr_decoded_andMatrixInput_1_8 }; 
    wire core_csr_decoded_andMatrixInput_7_6 = core_csr_decoded_plaInput_1 [29]; 
    wire core_csr_decoded_andMatrixInput_7_7 = core_csr_decoded_plaInput_1 [29]; 
    wire[1:0] core_csr_decoded_lo_lo_6 ={ core_csr_decoded_andMatrixInput_8_6 , core_csr_decoded_andMatrixInput_9_6 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_6 ={ core_csr_decoded_andMatrixInput_5_6 , core_csr_decoded_andMatrixInput_6_6 }; 
    wire[2:0] core_csr_decoded_lo_hi_6 ={ core_csr_decoded_lo_hi_hi_6 , core_csr_decoded_andMatrixInput_7_6 }; 
    wire[4:0] core_csr_decoded_lo_8 ={ core_csr_decoded_lo_hi_6 , core_csr_decoded_lo_lo_6 }; 
    wire[1:0] core_csr_decoded_hi_lo_6 ={ core_csr_decoded_andMatrixInput_3_8 , core_csr_decoded_andMatrixInput_4_6 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_6 ={ core_csr_decoded_andMatrixInput_0_9 , core_csr_decoded_andMatrixInput_1_9 }; 
    wire[2:0] core_csr_decoded_hi_hi_6 ={ core_csr_decoded_hi_hi_hi_6 , core_csr_decoded_andMatrixInput_2_8 }; 
    wire[4:0] core_csr_decoded_hi_8 ={ core_csr_decoded_hi_hi_6 , core_csr_decoded_hi_lo_6 }; 
    wire core_csr_decoded_andMatrixInput_0_10 = core_csr_decoded_plaInput_1 [22]; 
    wire[1:0] core_csr_decoded_lo_lo_7 ={ core_csr_decoded_andMatrixInput_8_7 , core_csr_decoded_andMatrixInput_9_7 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_7 ={ core_csr_decoded_andMatrixInput_5_7 , core_csr_decoded_andMatrixInput_6_7 }; 
    wire[2:0] core_csr_decoded_lo_hi_7 ={ core_csr_decoded_lo_hi_hi_7 , core_csr_decoded_andMatrixInput_7_7 }; 
    wire[4:0] core_csr_decoded_lo_9 ={ core_csr_decoded_lo_hi_7 , core_csr_decoded_lo_lo_7 }; 
    wire[1:0] core_csr_decoded_hi_lo_7 ={ core_csr_decoded_andMatrixInput_3_9 , core_csr_decoded_andMatrixInput_4_7 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_7 ={ core_csr_decoded_andMatrixInput_0_10 , core_csr_decoded_andMatrixInput_1_10 }; 
    wire[2:0] core_csr_decoded_hi_hi_7 ={ core_csr_decoded_hi_hi_hi_7 , core_csr_decoded_andMatrixInput_2_9 }; 
    wire[4:0] core_csr_decoded_hi_9 ={ core_csr_decoded_hi_hi_7 , core_csr_decoded_hi_lo_7 }; 
    wire core_csr_decoded_andMatrixInput_0_11 = core_csr_decoded_plaInput_1 [30]; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_lo_1 ={&{ core_csr_decoded_hi_9 , core_csr_decoded_lo_9 },&{ core_csr_decoded_hi_7 , core_csr_decoded_lo_7 }}; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_hi_hi_1 ={&{ core_csr_decoded_hi_5 , core_csr_decoded_lo_5 },&{ core_csr_decoded_hi_6 , core_csr_decoded_lo_6 }}; 
    wire[2:0] core_csr_decoded_orMatrixOutputs_hi_hi_1 ={ core_csr_decoded_orMatrixOutputs_hi_hi_hi_1 ,|{&{ core_csr_decoded_hi_8 , core_csr_decoded_lo_8 },&{ core_csr_decoded_andMatrixInput_0_11 , core_csr_decoded_andMatrixInput_1_11 }}}; 
    wire[4:0] core_csr_decoded_orMatrixOutputs_hi_1 ={ core_csr_decoded_orMatrixOutputs_hi_hi_1 , core_csr_decoded_orMatrixOutputs_hi_lo_1 }; 
    wire[8:0] core_csr_decoded_orMatrixOutputs_1 ={ core_csr_decoded_orMatrixOutputs_hi_1 ,4'h0}; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_lo_1 = core_csr_decoded_orMatrixOutputs_1 [1:0]; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_hi_1 = core_csr_decoded_orMatrixOutputs_1 [3:2]; 
    wire[3:0] core_csr_decoded_invMatrixOutputs_lo_1 ={ core_csr_decoded_invMatrixOutputs_lo_hi_1 , core_csr_decoded_invMatrixOutputs_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_lo_1 = core_csr_decoded_orMatrixOutputs_1 [5:4]; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_hi_hi_1 = core_csr_decoded_orMatrixOutputs_1 [8:7]; 
    wire[2:0] core_csr_decoded_invMatrixOutputs_hi_hi_1 ={ core_csr_decoded_invMatrixOutputs_hi_hi_hi_1 , core_csr_decoded_orMatrixOutputs_1 [6]}; 
    wire[4:0] core_csr_decoded_invMatrixOutputs_hi_1 ={ core_csr_decoded_invMatrixOutputs_hi_hi_1 , core_csr_decoded_invMatrixOutputs_hi_lo_1 }; 
  assign  core_csr_decoded_invMatrixOutputs_1 ={ core_csr_decoded_invMatrixOutputs_hi_1 , core_csr_decoded_invMatrixOutputs_lo_1 }; 
    wire[8:0] core_csr_decoded_196 = core_csr_decoded_invMatrixOutputs_1 ; 
    wire core_csr_is_break = core_csr_decoded_196 [7]; 
    wire core_csr_is_ret = core_csr_decoded_196 [6]; 
    wire core_csr_is_wfi = core_csr_decoded_196 [4]; 
    wire core_csr_is_sfence = core_csr_decoded_196 [3]; 
    wire core_csr_is_hfence_vvma = core_csr_decoded_196 [2]; 
    wire core_csr_is_hfence_gvma = core_csr_decoded_196 [1]; 
    wire core_csr_is_hlsv = core_csr_decoded_196 [0]; 
    wire core_csr_is_counter = core_csr_addr_1 >12'hBFF& core_csr_addr_1 <12'hC20| core_csr_addr_1 >12'hC7F& core_csr_addr_1 <12'hCA0; 
    wire[4:0] core_csr_counter_addr = core_csr_addr_1 [4:0]; 
    wire[31:0] core_csr__GEN_4 ={27'h0, core_csr_counter_addr }; 
    wire[31:0] core_csr__io_decode_0_virtual_access_illegal_T_3 =32'h0>> core_csr__GEN_4 ; 
    wire[31:0] core_csr__io_decode_0_virtual_access_illegal_T_6 =32'h0>> core_csr__GEN_4 ; 
    wire[11:0] core_csr_io_decode_0_fp_csr_invInputs =~ core_csr_io_decode_0_fp_csr_plaInput ; 
    wire core_csr_csr_exists = core_csr_addr_1 ==12'h7A0| core_csr_addr_1 ==12'h7A1| core_csr_addr_1 ==12'h7A2| core_csr_addr_1 ==12'h7A3| core_csr_addr_1 ==12'h301| core_csr_addr_1 ==12'h300| core_csr_addr_1 ==12'h305| core_csr_addr_1 ==12'h344| core_csr_addr_1 ==12'h304| core_csr_addr_1 ==12'h340| core_csr_addr_1 ==12'h341| core_csr_addr_1 ==12'h343| core_csr_addr_1 ==12'h342| core_csr_addr_1 ==12'hF14| core_csr_addr_1 ==12'h7B0| core_csr_addr_1 ==12'h7B1| core_csr_addr_1 ==12'h7B2| core_csr_addr_1 ==12'h320| core_csr_addr_1 ==12'hB00| core_csr_addr_1 ==12'hB02| core_csr_addr_1 ==12'h323| core_csr_addr_1 ==12'hB03| core_csr_addr_1 ==12'hC03| core_csr_addr_1 ==12'hB83| core_csr_addr_1 ==12'hC83| core_csr_addr_1 ==12'h324| core_csr_addr_1 ==12'hB04| core_csr_addr_1 ==12'hC04| core_csr_addr_1 ==12'hB84| core_csr_addr_1 ==12'hC84| core_csr_addr_1 ==12'h325| core_csr_addr_1 ==12'hB05| core_csr_addr_1 ==12'hC05| core_csr_addr_1 ==12'hB85| core_csr_addr_1 ==12'hC85| core_csr_addr_1 ==12'h326| core_csr_addr_1 ==12'hB06| core_csr_addr_1 ==12'hC06| core_csr_addr_1 ==12'hB86| core_csr_addr_1 ==12'hC86| core_csr_addr_1 ==12'h327| core_csr_addr_1 ==12'hB07| core_csr_addr_1 ==12'hC07| core_csr_addr_1 ==12'hB87| core_csr_addr_1 ==12'hC87| core_csr_addr_1 ==12'h328| core_csr_addr_1 ==12'hB08| core_csr_addr_1 ==12'hC08| core_csr_addr_1 ==12'hB88| core_csr_addr_1 ==12'hC88| core_csr_addr_1 ==12'h329| core_csr_addr_1 ==12'hB09| core_csr_addr_1 ==12'hC09| core_csr_addr_1 ==12'hB89| core_csr_addr_1 ==12'hC89| core_csr_addr_1 ==12'h32A| core_csr_addr_1 ==12'hB0A| core_csr_addr_1 ==12'hC0A| core_csr_addr_1 ==12'hB8A| core_csr_addr_1 ==12'hC8A| core_csr_addr_1 ==12'h32B| core_csr_addr_1 ==12'hB0B| core_csr_addr_1 ==12'hC0B| core_csr_addr_1 ==12'hB8B| core_csr_addr_1 ==12'hC8B| core_csr_addr_1 ==12'h32C| core_csr_addr_1 ==12'hB0C| core_csr_addr_1 ==12'hC0C| core_csr_addr_1 ==12'hB8C| core_csr_addr_1 ==12'hC8C| core_csr_addr_1 ==12'h32D| core_csr_addr_1 ==12'hB0D| core_csr_addr_1 ==12'hC0D| core_csr_addr_1 ==12'hB8D| core_csr_addr_1 ==12'hC8D| core_csr_addr_1 ==12'h32E| core_csr_addr_1 ==12'hB0E| core_csr_addr_1 ==12'hC0E| core_csr_addr_1 ==12'hB8E| core_csr_addr_1 ==12'hC8E| core_csr_addr_1 ==12'h32F| core_csr_addr_1 ==12'hB0F| core_csr_addr_1 ==12'hC0F| core_csr_addr_1 ==12'hB8F| core_csr_addr_1 ==12'hC8F| core_csr_addr_1 ==12'h330| core_csr_addr_1 ==12'hB10| core_csr_addr_1 ==12'hC10| core_csr_addr_1 ==12'hB90| core_csr_addr_1 ==12'hC90| core_csr_addr_1 ==12'h331| core_csr_addr_1 ==12'hB11| core_csr_addr_1 ==12'hC11| core_csr_addr_1 ==12'hB91| core_csr_addr_1 ==12'hC91| core_csr_addr_1 ==12'h332| core_csr_addr_1 ==12'hB12| core_csr_addr_1 ==12'hC12| core_csr_addr_1 ==12'hB92| core_csr_addr_1 ==12'hC92| core_csr_addr_1 ==12'h333| core_csr_addr_1 ==12'hB13| core_csr_addr_1 ==12'hC13| core_csr_addr_1 ==12'hB93| core_csr_addr_1 ==12'hC93| core_csr_addr_1 ==12'h334| core_csr_addr_1 ==12'hB14| core_csr_addr_1 ==12'hC14| core_csr_addr_1 ==12'hB94| core_csr_addr_1 ==12'hC94| core_csr_addr_1 ==12'h335| core_csr_addr_1 ==12'hB15| core_csr_addr_1 ==12'hC15| core_csr_addr_1 ==12'hB95| core_csr_addr_1 ==12'hC95| core_csr_addr_1 ==12'h336| core_csr_addr_1 ==12'hB16| core_csr_addr_1 ==12'hC16| core_csr_addr_1 ==12'hB96| core_csr_addr_1 ==12'hC96| core_csr_addr_1 ==12'h337| core_csr_addr_1 ==12'hB17| core_csr_addr_1 ==12'hC17| core_csr_addr_1 ==12'hB97| core_csr_addr_1 ==12'hC97| core_csr_addr_1 ==12'h338| core_csr_addr_1 ==12'hB18| core_csr_addr_1 ==12'hC18| core_csr_addr_1 ==12'hB98| core_csr_addr_1 ==12'hC98| core_csr_addr_1 ==12'h339| core_csr_addr_1 ==12'hB19| core_csr_addr_1 ==12'hC19| core_csr_addr_1 ==12'hB99| core_csr_addr_1 ==12'hC99| core_csr_addr_1 ==12'h33A| core_csr_addr_1 ==12'hB1A| core_csr_addr_1 ==12'hC1A| core_csr_addr_1 ==12'hB9A| core_csr_addr_1 ==12'hC9A| core_csr_addr_1 ==12'h33B| core_csr_addr_1 ==12'hB1B| core_csr_addr_1 ==12'hC1B| core_csr_addr_1 ==12'hB9B| core_csr_addr_1 ==12'hC9B| core_csr_addr_1 ==12'h33C| core_csr_addr_1 ==12'hB1C| core_csr_addr_1 ==12'hC1C| core_csr_addr_1 ==12'hB9C| core_csr_addr_1 ==12'hC9C| core_csr_addr_1 ==12'h33D| core_csr_addr_1 ==12'hB1D| core_csr_addr_1 ==12'hC1D| core_csr_addr_1 ==12'hB9D| core_csr_addr_1 ==12'hC9D| core_csr_addr_1 ==12'h33E| core_csr_addr_1 ==12'hB1E| core_csr_addr_1 ==12'hC1E| core_csr_addr_1 ==12'hB9E| core_csr_addr_1 ==12'hC9E| core_csr_addr_1 ==12'h33F| core_csr_addr_1 ==12'hB1F| core_csr_addr_1 ==12'hC1F| core_csr_addr_1 ==12'hB9F| core_csr_addr_1 ==12'hC9F| core_csr_addr_1 ==12'hC00| core_csr_addr_1 ==12'hC02| core_csr_addr_1 ==12'hB80| core_csr_addr_1 ==12'hB82| core_csr_addr_1 ==12'hC80| core_csr_addr_1 ==12'hC82| core_csr_addr_1 ==12'h3A0| core_csr_addr_1 ==12'h3A1| core_csr_addr_1 ==12'h3A2| core_csr_addr_1 ==12'h3A3| core_csr_addr_1 ==12'h3B0| core_csr_addr_1 ==12'h3B1| core_csr_addr_1 ==12'h3B2| core_csr_addr_1 ==12'h3B3| core_csr_addr_1 ==12'h3B4| core_csr_addr_1 ==12'h3B5| core_csr_addr_1 ==12'h3B6| core_csr_addr_1 ==12'h3B7| core_csr_addr_1 ==12'h3B8| core_csr_addr_1 ==12'h3B9| core_csr_addr_1 ==12'h3BA| core_csr_addr_1 ==12'h3BB| core_csr_addr_1 ==12'h3BC| core_csr_addr_1 ==12'h3BD| core_csr_addr_1 ==12'h3BE| core_csr_addr_1 ==12'h3BF| core_csr_addr_1 ==12'h7C1| core_csr_addr_1 ==12'hF12| core_csr_addr_1 ==12'hF11| core_csr_addr_1 ==12'hF13| core_csr_addr_1 ==12'hF15; 
    wire[11:0] core_csr_io_decode_0_read_illegal_invInputs =~ core_csr_io_decode_0_read_illegal_plaInput ; 
    wire core_csr_io_decode_0_read_illegal_invMatrixOutputs ; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_0 = core_csr_io_decode_0_read_illegal_plaInput [4]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_1 = core_csr_io_decode_0_read_illegal_plaInput [5]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_2 = core_csr_io_decode_0_read_illegal_invInputs [6]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_3 = core_csr_io_decode_0_read_illegal_plaInput [7]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_4 = core_csr_io_decode_0_read_illegal_plaInput [8]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_5 = core_csr_io_decode_0_read_illegal_plaInput [9]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_6 = core_csr_io_decode_0_read_illegal_plaInput [10]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_7 = core_csr_io_decode_0_read_illegal_invInputs [11]; 
    wire[1:0] core_csr_io_decode_0_read_illegal_lo_lo ={ core_csr_io_decode_0_read_illegal_andMatrixInput_6 , core_csr_io_decode_0_read_illegal_andMatrixInput_7 }; 
    wire[1:0] core_csr_io_decode_0_read_illegal_lo_hi ={ core_csr_io_decode_0_read_illegal_andMatrixInput_4 , core_csr_io_decode_0_read_illegal_andMatrixInput_5 }; 
    wire[3:0] core_csr_io_decode_0_read_illegal_lo ={ core_csr_io_decode_0_read_illegal_lo_hi , core_csr_io_decode_0_read_illegal_lo_lo }; 
    wire[1:0] core_csr_io_decode_0_read_illegal_hi_lo ={ core_csr_io_decode_0_read_illegal_andMatrixInput_2 , core_csr_io_decode_0_read_illegal_andMatrixInput_3 }; 
    wire[1:0] core_csr_io_decode_0_read_illegal_hi_hi ={ core_csr_io_decode_0_read_illegal_andMatrixInput_0 , core_csr_io_decode_0_read_illegal_andMatrixInput_1 }; 
    wire[3:0] core_csr_io_decode_0_read_illegal_hi ={ core_csr_io_decode_0_read_illegal_hi_hi , core_csr_io_decode_0_read_illegal_hi_lo }; 
    wire core_csr_io_decode_0_read_illegal_orMatrixOutputs =&{ core_csr_io_decode_0_read_illegal_hi , core_csr_io_decode_0_read_illegal_lo }; 
  assign  core_csr_io_decode_0_read_illegal_invMatrixOutputs = core_csr_io_decode_0_read_illegal_orMatrixOutputs ; 
    wire core_csr_io_decode_0_read_illegal_plaOutput = core_csr_io_decode_0_read_illegal_invMatrixOutputs ; 
    wire[11:0] core_csr_io_decode_0_read_illegal_invInputs_1 =~ core_csr_io_decode_0_read_illegal_plaInput_1 ; 
    wire[11:0] core_csr_io_decode_0_write_flush_addr_m ={ core_csr_addr_1 [11:10], core_csr_addr_1 [9:0]|10'h300}; 
    wire[31:0] core_csr_cause = core_csr_insn_call  ? {28'h0,{3'h1,~ core_csr_reg_mstatus_v }-4'h8}: core_csr_insn_break  ? 32'h3: core_csr_io_cause ; 
    wire[7:0] core_csr_cause_lsbs = core_csr_cause [7:0]; 
    wire core_csr__causeIsDebugTrigger_T_2 = core_csr_cause_lsbs ==8'hE; 
    wire core_csr_causeIsDebugInt = core_csr_cause [31]& core_csr__causeIsDebugTrigger_T_2 ; 
    wire core_csr_causeIsDebugTrigger =~( core_csr_cause [31])& core_csr__causeIsDebugTrigger_T_2 ; 
    wire[1:0] core_csr_causeIsDebugBreak_hi ={ core_csr_reg_dcsr_ebreakm ,1'h0}; 
    wire core_csr_causeIsDebugBreak =~( core_csr_cause [31])& core_csr_insn_break & core_csr_causeIsDebugBreak_hi [1]; 
    wire core_csr_trapToDebug = core_csr_reg_singleStepped | core_csr_causeIsDebugInt | core_csr_causeIsDebugTrigger | core_csr_causeIsDebugBreak | core_csr_reg_debug ; 
    wire[11:0] core_csr_debugTVec = core_csr_reg_debug  ? {8'h80,~ core_csr_insn_break ,3'h0}:12'h800; 
    wire[6:0] core_csr_notDebugTVec_interruptOffset ={ core_csr_cause [4:0],2'h0}; 
    wire[31:0] core_csr_notDebugTVec_interruptVec ={ core_csr_notDebugTVec_base [31:7], core_csr_notDebugTVec_interruptOffset }; 
    wire core_csr_notDebugTVec_doVector = core_csr_notDebugTVec_base [0]& core_csr_cause [31]& core_csr_cause_lsbs [7:5]==3'h0; 
    wire[31:0] core_csr_notDebugTVec = core_csr_notDebugTVec_doVector  ?  core_csr_notDebugTVec_interruptVec :{ core_csr_notDebugTVec_base [31:2],2'h0}; 
    wire core_csr__causeIsRnmiBEU_T_3 = core_csr_cause_lsbs ==8'hC; 
    wire core_csr_causeIsRnmiInt = core_csr_cause [31]& core_csr_cause [30]&( core_csr_cause_lsbs ==8'hD| core_csr__causeIsRnmiBEU_T_3 ); 
    wire core_csr_causeIsRnmiBEU = core_csr_cause [31]& core_csr_cause [30]& core_csr__causeIsRnmiBEU_T_3 ; 
    wire[31:0] core_csr_tvec = core_csr_trapToDebug  ? {20'h0, core_csr_debugTVec }: core_csr_notDebugTVec ; 
    wire core_csr__exception_T = core_csr_insn_call | core_csr_insn_break ; 
  assign  core_csr__io_singleStep_output = core_csr_reg_dcsr_step &~ core_csr_reg_debug ; 
    wire core_csr_exception = core_csr__exception_T | core_csr_io_exception ; 
    wire[2:0] core_csr__GEN_5 ={1'h0,{1'h0, core_csr_insn_ret }+{1'h0, core_csr_insn_call }}+{1'h0,{1'h0, core_csr_insn_break }+{1'h0, core_csr_io_exception }}; 
  always @( posedge  core_csr_clock )
         begin 
             if (~ core_csr_reset &(|( core_csr__GEN_5 [2:1])))
                 begin 
                     if (1)$error("Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:1010 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1.U, \"these conditions must be mutually exclusive\")\n");
                     if (1)$fatal;
                 end 
             if (~ core_csr_reset &~(~ core_csr_reg_singleStepped |~ core_csr_io_retire ))
                 begin 
                     if (1)$error("Assertion failed\n    at CSR.scala:1019 assert(!reg_singleStepped || io.retire === 0.U)\n");
                     if (1)$fatal;
                 end 
         end
    wire[31:0] core_csr_epc ={ core_csr_io_pc [31:1],1'h0}; 
    wire[31:0] core_csr_tval = core_csr_insn_break  ?  core_csr_epc : core_csr_io_tval ; 
    wire core_csr_en_3 = core_csr_exception & core_csr_cause ==32'h80000003; 
    wire core_csr_en_7 = core_csr_exception & core_csr_cause ==32'h80000007; 
    wire core_csr_en_11 = core_csr_exception & core_csr_cause ==32'h8000000B; 
    wire core_csr_en_16 = core_csr_exception & core_csr_cause ==32'h0; 
    wire core_csr_en_17 = core_csr_exception & core_csr_cause ==32'h1; 
    wire core_csr_en_18 = core_csr_exception & core_csr_cause ==32'h2; 
    wire core_csr_en_19 = core_csr_exception & core_csr_cause ==32'h3; 
    wire core_csr_en_20 = core_csr_exception & core_csr_cause ==32'h4; 
    wire core_csr_en_21 = core_csr_exception & core_csr_cause ==32'h5; 
    wire core_csr_en_22 = core_csr_exception & core_csr_cause ==32'h6; 
    wire core_csr_en_23 = core_csr_exception & core_csr_cause ==32'h7; 
    wire core_csr_en_24 = core_csr_exception & core_csr_cause ==32'hB; 
    wire core_csr__GEN_6 = core_csr_io_rw_addr [10]& core_csr_io_rw_addr [7]; 
    wire[1:0] core_csr_ret_prv = core_csr__GEN_6  ? 2'h3: core_csr_reg_mstatus_mpp ; 
    wire[1:0] core_csr_new_prv = core_csr_insn_ret  ?  core_csr_ret_prv :2'h3; 
  assign  core_csr__io_csr_stall_output = core_csr_reg_wfi | core_csr_io_status_cease_r ; 
    wire[31:0] core_csr__io_rw_rdata_T_197 =( core_csr_decoded_1  ? { core_csr_hi_4 , core_csr_lo_4 }:32'h0)|( core_csr_decoded_2  ?  core_csr_reg_bp_0_address :32'h0); 
    wire[31:0] core_csr__io_rw_rdata_T_201 ={ core_csr__io_rw_rdata_T_197 [31:26], core_csr__io_rw_rdata_T_197 [25:0]|( core_csr_decoded_3  ? { core_csr_hi_5 , core_csr_lo_5 }:26'h0)}|( core_csr_decoded_4  ?  core_csr_reg_misa :32'h0)|( core_csr_decoded_5  ?  core_csr_read_mstatus :32'h0)|( core_csr_decoded_6  ?  core_csr_read_mtvec :32'h0); 
    wire[31:0] core_csr__io_rw_rdata_T_207 ={ core_csr__io_rw_rdata_T_201 [31:16], core_csr__io_rw_rdata_T_201 [15:0]|( core_csr_decoded_7  ?  core_csr_read_mip :16'h0)}|( core_csr_decoded_8  ?  core_csr_reg_mie :32'h0)|( core_csr_decoded_9  ?  core_csr_reg_mscratch :32'h0)|( core_csr_decoded_10  ? ~{ core_csr__io_evec_T_20 [31:2], core_csr__io_evec_T_20 [1:0]| core_csr__GEN_3 }:32'h0)|( core_csr_decoded_11  ?  core_csr_reg_mtval :32'h0)|( core_csr_decoded_12  ?  core_csr_reg_mcause :32'h0); 
    wire[31:0] core_csr__io_rw_rdata_T_211 ={ core_csr__io_rw_rdata_T_207 [31:1], core_csr__io_rw_rdata_T_207 [0]| core_csr_decoded_13 & core_csr_io_hartid }|( core_csr_decoded_14  ? { core_csr_hi_6 , core_csr_lo_6 }:32'h0)|( core_csr_decoded_15  ? ~{ core_csr__io_evec_T_10 [31:2], core_csr__io_evec_T_10 [1:0]| core_csr__GEN_3 }:32'h0)|( core_csr_decoded_16  ?  core_csr_reg_dscratch0 :32'h0); 
    wire[31:0] core_csr__GEN_7 ={ core_csr__io_rw_rdata_T_211 [31:3], core_csr__io_rw_rdata_T_211 [2:0]|( core_csr_decoded_17  ?  core_csr_reg_mcountinhibit :3'h0)}|( core_csr_decoded_18  ?  core_csr_value_1 [31:0]:32'h0)|( core_csr_decoded_19  ?  core_csr_value [31:0]:32'h0)|( core_csr_decoded_165  ?  core_csr_value_1 [31:0]:32'h0)|( core_csr_decoded_166  ?  core_csr_value [31:0]:32'h0)|( core_csr_decoded_167  ?  core_csr_value_1 [63:32]:32'h0)|( core_csr_decoded_168  ?  core_csr_value [63:32]:32'h0)|( core_csr_decoded_169  ?  core_csr_value_1 [63:32]:32'h0)|( core_csr_decoded_170  ?  core_csr_value [63:32]:32'h0)|( core_csr_decoded_171  ? { core_csr_hi_11 , core_csr_lo_11 }:32'h0)|( core_csr_decoded_172  ? { core_csr_hi_16 , core_csr_lo_16 }:32'h0); 
    wire[29:0] core_csr__GEN_8 = core_csr__GEN_7 [29:0]|( core_csr_decoded_175  ?  core_csr_reg_pmp_0_addr :30'h0)|( core_csr_decoded_176  ?  core_csr_reg_pmp_1_addr :30'h0)|( core_csr_decoded_177  ?  core_csr_reg_pmp_2_addr :30'h0)|( core_csr_decoded_178  ?  core_csr_reg_pmp_3_addr :30'h0)|( core_csr_decoded_179  ?  core_csr_reg_pmp_4_addr :30'h0)|( core_csr_decoded_180  ?  core_csr_reg_pmp_5_addr :30'h0)|( core_csr_decoded_181  ?  core_csr_reg_pmp_6_addr :30'h0)|( core_csr_decoded_182  ?  core_csr_reg_pmp_7_addr :30'h0); 
  assign  core_csr__io_rw_rdata_output =( core_csr_decoded_191  ?  core_csr_reg_custom_0 :32'h0)|{ core_csr__GEN_7 [31:30], core_csr__GEN_8 [29:1], core_csr__GEN_8 [0]| core_csr_decoded_192 }|( core_csr_decoded_194  ? 32'h20181004:32'h0); 
    wire core_csr_csr_wen = core_csr_io_rw_cmd ==3'h6|(& core_csr_io_rw_cmd )| core_csr_io_rw_cmd ==3'h5; 
    wire core_csr_new_mstatus_uie = core_csr_wdata [0]; 
    wire core_csr_new_mstatus_sie = core_csr_wdata [1]; 
    wire core_csr_new_mstatus_hie = core_csr_wdata [2]; 
    wire core_csr_new_mstatus_mie = core_csr_wdata [3]; 
    wire core_csr_new_mstatus_upie = core_csr_wdata [4]; 
    wire core_csr_new_mstatus_spie = core_csr_wdata [5]; 
    wire core_csr_new_mstatus_ube = core_csr_wdata [6]; 
    wire core_csr_new_mstatus_mpie = core_csr_wdata [7]; 
    wire core_csr_new_mstatus_spp = core_csr_wdata [8]; 
    wire[1:0] core_csr_new_mstatus_vs = core_csr_wdata [10:9]; 
    wire[1:0] core_csr_new_mstatus_mpp = core_csr_wdata [12:11]; 
    wire[1:0] core_csr_new_mstatus_fs = core_csr_wdata [14:13]; 
    wire[1:0] core_csr_new_mstatus_xs = core_csr_wdata [16:15]; 
    wire core_csr_new_mstatus_mprv = core_csr_wdata [17]; 
    wire core_csr_new_mstatus_sum = core_csr_wdata [18]; 
    wire core_csr_new_mstatus_mxr = core_csr_wdata [19]; 
    wire core_csr_new_mstatus_tvm = core_csr_wdata [20]; 
    wire core_csr_new_mstatus_tw = core_csr_wdata [21]; 
    wire core_csr_new_mstatus_tsr = core_csr_wdata [22]; 
    wire[7:0] core_csr_new_mstatus_zero1 = core_csr_wdata [30:23]; 
    wire core_csr_new_mstatus_sd_rv32 = core_csr_wdata [31]; 
    wire core_csr_f = core_csr_wdata [5]; 
    wire[3:0] core_csr_new_mip_lo_lo ={ core_csr_new_mip_lo_lo_hi , core_csr_new_mip_lo_lo_lo }; 
    wire[3:0] core_csr_new_mip_lo_hi ={ core_csr_new_mip_lo_hi_hi , core_csr_new_mip_lo_hi_lo }; 
    wire[7:0] core_csr_new_mip_lo ={ core_csr_new_mip_lo_hi , core_csr_new_mip_lo_lo }; 
    wire[3:0] core_csr_new_mip_hi_lo ={ core_csr_new_mip_hi_lo_hi , core_csr_new_mip_hi_lo_lo }; 
    wire[3:0] core_csr_new_mip_hi_hi ={ core_csr_new_mip_hi_hi_hi , core_csr_new_mip_hi_hi_lo }; 
    wire[7:0] core_csr_new_mip_hi ={ core_csr_new_mip_hi_hi , core_csr_new_mip_hi_lo }; 
    wire[15:0] core_csr__new_mip_WIRE =(( core_csr_io_rw_cmd [1] ? { core_csr_new_mip_hi , core_csr_new_mip_lo }:16'h0)| core_csr_io_rw_wdata [15:0])&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata [15:0]:16'h0); 
    wire core_csr_new_mip_usip = core_csr__new_mip_WIRE [0]; 
    wire core_csr_new_mip_ssip = core_csr__new_mip_WIRE [1]; 
    wire core_csr_new_mip_vssip = core_csr__new_mip_WIRE [2]; 
    wire core_csr_new_mip_msip = core_csr__new_mip_WIRE [3]; 
    wire core_csr_new_mip_utip = core_csr__new_mip_WIRE [4]; 
    wire core_csr_new_mip_stip = core_csr__new_mip_WIRE [5]; 
    wire core_csr_new_mip_vstip = core_csr__new_mip_WIRE [6]; 
    wire core_csr_new_mip_mtip = core_csr__new_mip_WIRE [7]; 
    wire core_csr_new_mip_ueip = core_csr__new_mip_WIRE [8]; 
    wire core_csr_new_mip_seip = core_csr__new_mip_WIRE [9]; 
    wire core_csr_new_mip_vseip = core_csr__new_mip_WIRE [10]; 
    wire core_csr_new_mip_meip = core_csr__new_mip_WIRE [11]; 
    wire core_csr_new_mip_sgeip = core_csr__new_mip_WIRE [12]; 
    wire core_csr_new_mip_rocc = core_csr__new_mip_WIRE [13]; 
    wire core_csr_new_mip_debug = core_csr__new_mip_WIRE [14]; 
    wire core_csr_new_mip_zero1 = core_csr__new_mip_WIRE [15]; 
    wire[1:0] core_csr_new_dcsr_prv = core_csr_wdata [1:0]; 
    wire core_csr_new_dcsr_step = core_csr_wdata [2]; 
    wire[1:0] core_csr_new_dcsr_zero1 = core_csr_wdata [4:3]; 
    wire core_csr_new_dcsr_v = core_csr_wdata [5]; 
    wire[2:0] core_csr_new_dcsr_cause = core_csr_wdata [8:6]; 
    wire core_csr_new_dcsr_stoptime = core_csr_wdata [9]; 
    wire core_csr_new_dcsr_stopcycle = core_csr_wdata [10]; 
    wire core_csr_new_dcsr_zero2 = core_csr_wdata [11]; 
    wire core_csr_new_dcsr_ebreaku = core_csr_wdata [12]; 
    wire core_csr_new_dcsr_ebreaks = core_csr_wdata [13]; 
    wire core_csr_new_dcsr_ebreakh = core_csr_wdata [14]; 
    wire core_csr_new_dcsr_ebreakm = core_csr_wdata [15]; 
    wire[11:0] core_csr_new_dcsr_zero3 = core_csr_wdata [27:16]; 
    wire[1:0] core_csr_new_dcsr_zero4 = core_csr_wdata [29:28]; 
    wire[1:0] core_csr_new_dcsr_xdebugver = core_csr_wdata [31:30]; 
    wire[2:0] core_csr_newBPC_lo_lo ={ core_csr_newBPC_lo_lo_hi , core_csr_reg_bp_0_control_r }; 
    wire[6:0] core_csr_newBPC_lo ={4'h8, core_csr_newBPC_lo_lo }; 
    wire[5:0] core_csr_newBPC_hi_lo ={ core_csr_newBPC_hi_lo_hi , core_csr_newBPC_hi_lo_lo }; 
    wire[18:0] core_csr_newBPC_hi_hi ={ core_csr_newBPC_hi_hi_hi ,14'h400}; 
    wire[24:0] core_csr_newBPC_hi ={ core_csr_newBPC_hi_hi , core_csr_newBPC_hi_lo }; 
    wire[31:0] core_csr__newBPC_WIRE =(( core_csr_io_rw_cmd [1] ? { core_csr_newBPC_hi , core_csr_newBPC_lo }:32'h0)| core_csr_io_rw_wdata )&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :32'h0); 
    wire core_csr_newBPC_r = core_csr__newBPC_WIRE [0]; 
    wire core_csr_newBPC_w = core_csr__newBPC_WIRE [1]; 
    wire core_csr_newBPC_x = core_csr__newBPC_WIRE [2]; 
    wire core_csr_newBPC_u = core_csr__newBPC_WIRE [3]; 
    wire core_csr_newBPC_s = core_csr__newBPC_WIRE [4]; 
    wire core_csr_newBPC_h = core_csr__newBPC_WIRE [5]; 
    wire core_csr_newBPC_m = core_csr__newBPC_WIRE [6]; 
    wire[1:0] core_csr_newBPC_tmatch = core_csr__newBPC_WIRE [8:7]; 
    wire[1:0] core_csr_newBPC_zero = core_csr__newBPC_WIRE [10:9]; 
    wire core_csr_newBPC_chain = core_csr__newBPC_WIRE [11]; 
    wire core_csr_newBPC_action = core_csr__newBPC_WIRE [12]; 
    wire[7:0] core_csr_newBPC_reserved = core_csr__newBPC_WIRE [20:13]; 
    wire[5:0] core_csr_newBPC_maskmax = core_csr__newBPC_WIRE [26:21]; 
    wire core_csr_newBPC_dmode = core_csr__newBPC_WIRE [27]; 
    wire[3:0] core_csr_newBPC_ttype = core_csr__newBPC_WIRE [31:28]; 
    wire core_csr_dMode = core_csr_newBPC_dmode & core_csr_reg_debug ; 
    wire[31:0] core_csr__newBPC_WIRE_1 = core_csr_io_rw_wdata &~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :32'h0); 
    wire core_csr_newBPC_1_r = core_csr__newBPC_WIRE_1 [0]; 
    wire core_csr_newBPC_1_w = core_csr__newBPC_WIRE_1 [1]; 
    wire core_csr_newBPC_1_x = core_csr__newBPC_WIRE_1 [2]; 
    wire core_csr_newBPC_1_u = core_csr__newBPC_WIRE_1 [3]; 
    wire core_csr_newBPC_1_s = core_csr__newBPC_WIRE_1 [4]; 
    wire core_csr_newBPC_1_h = core_csr__newBPC_WIRE_1 [5]; 
    wire core_csr_newBPC_1_m = core_csr__newBPC_WIRE_1 [6]; 
    wire[1:0] core_csr_newBPC_1_tmatch = core_csr__newBPC_WIRE_1 [8:7]; 
    wire[1:0] core_csr_newBPC_1_zero = core_csr__newBPC_WIRE_1 [10:9]; 
    wire core_csr_newBPC_1_chain = core_csr__newBPC_WIRE_1 [11]; 
    wire core_csr_newBPC_1_action = core_csr__newBPC_WIRE_1 [12]; 
    wire[7:0] core_csr_newBPC_1_reserved = core_csr__newBPC_WIRE_1 [20:13]; 
    wire[5:0] core_csr_newBPC_1_maskmax = core_csr__newBPC_WIRE_1 [26:21]; 
    wire core_csr_newBPC_1_dmode = core_csr__newBPC_WIRE_1 [27]; 
    wire[3:0] core_csr_newBPC_1_ttype = core_csr__newBPC_WIRE_1 [31:28]; 
    wire core_csr_dMode_1 = core_csr_newBPC_1_dmode & core_csr_reg_debug ; 
    wire core_csr_newCfg_r = core_csr_wdata [0]; 
    wire core_csr_newCfg_w = core_csr_wdata [1]; 
    wire core_csr_newCfg_x = core_csr_wdata [2]; 
    wire[1:0] core_csr_newCfg_a = core_csr_wdata [4:3]; 
    wire[1:0] core_csr_newCfg_res = core_csr_wdata [6:5]; 
    wire core_csr_newCfg_l = core_csr_wdata [7]; 
    wire core_csr_newCfg_1_r = core_csr_wdata [8]; 
    wire core_csr_newCfg_1_w = core_csr_wdata [9]; 
    wire core_csr_newCfg_1_x = core_csr_wdata [10]; 
    wire[1:0] core_csr_newCfg_1_a = core_csr_wdata [12:11]; 
    wire[1:0] core_csr_newCfg_1_res = core_csr_wdata [14:13]; 
    wire core_csr_newCfg_1_l = core_csr_wdata [15]; 
    wire core_csr_newCfg_2_r = core_csr_wdata [16]; 
    wire core_csr_newCfg_2_w = core_csr_wdata [17]; 
    wire core_csr_newCfg_2_x = core_csr_wdata [18]; 
    wire[1:0] core_csr_newCfg_2_a = core_csr_wdata [20:19]; 
    wire[1:0] core_csr_newCfg_2_res = core_csr_wdata [22:21]; 
    wire core_csr_newCfg_2_l = core_csr_wdata [23]; 
    wire core_csr_newCfg_3_r = core_csr_wdata [24]; 
    wire core_csr_newCfg_3_w = core_csr_wdata [25]; 
    wire core_csr_newCfg_3_x = core_csr_wdata [26]; 
    wire[1:0] core_csr_newCfg_3_a = core_csr_wdata [28:27]; 
    wire[1:0] core_csr_newCfg_3_res = core_csr_wdata [30:29]; 
    wire core_csr_newCfg_3_l = core_csr_wdata [31]; 
    wire core_csr_newCfg_4_r = core_csr_wdata [0]; 
    wire core_csr_newCfg_4_w = core_csr_wdata [1]; 
    wire core_csr_newCfg_4_x = core_csr_wdata [2]; 
    wire[1:0] core_csr_newCfg_4_a = core_csr_wdata [4:3]; 
    wire[1:0] core_csr_newCfg_4_res = core_csr_wdata [6:5]; 
    wire core_csr_newCfg_4_l = core_csr_wdata [7]; 
    wire core_csr_newCfg_5_r = core_csr_wdata [8]; 
    wire core_csr_newCfg_5_w = core_csr_wdata [9]; 
    wire core_csr_newCfg_5_x = core_csr_wdata [10]; 
    wire[1:0] core_csr_newCfg_5_a = core_csr_wdata [12:11]; 
    wire[1:0] core_csr_newCfg_5_res = core_csr_wdata [14:13]; 
    wire core_csr_newCfg_5_l = core_csr_wdata [15]; 
    wire core_csr_newCfg_6_r = core_csr_wdata [16]; 
    wire core_csr_newCfg_6_w = core_csr_wdata [17]; 
    wire core_csr_newCfg_6_x = core_csr_wdata [18]; 
    wire[1:0] core_csr_newCfg_6_a = core_csr_wdata [20:19]; 
    wire[1:0] core_csr_newCfg_6_res = core_csr_wdata [22:21]; 
    wire core_csr_newCfg_6_l = core_csr_wdata [23]; 
    wire core_csr_newCfg_7_r = core_csr_wdata [24]; 
    wire core_csr_newCfg_7_w = core_csr_wdata [25]; 
    wire core_csr_newCfg_7_x = core_csr_wdata [26]; 
    wire[1:0] core_csr_newCfg_7_a = core_csr_wdata [28:27]; 
    wire[1:0] core_csr_newCfg_7_res = core_csr_wdata [30:29]; 
    wire core_csr_newCfg_7_l = core_csr_wdata [31]; 
    wire[31:0] core_csr__reg_misa_T =~ core_csr_wdata ; 
    wire core_csr__large_T_2 = core_csr_nextSmall [6]&~ core_csr_x3 ; 
    wire[57:0] core_csr__large_r_T = core_csr_large_0 +58'h1; 
    wire core_csr__GEN_9 =~ core_csr_insn_ret | core_csr__GEN_6 ; 
    wire core_csr__GEN_10 = core_csr_exception & core_csr_trapToDebug &~ core_csr_reg_debug ; 
    wire core_csr__GEN_11 =~ core_csr_exception | core_csr_trapToDebug ; 
    wire core_csr__GEN_12 =~ core_csr_reg_bp_0_control_dmode | core_csr_reg_debug ; 
    wire core_csr__GEN_13 = core_csr_csr_wen & core_csr__GEN_12 & core_csr_decoded_1 ; 
    wire core_csr__GEN_14 = core_csr_csr_wen & core_csr_decoded_171 &~ core_csr_reg_pmp_0_cfg_l ; 
    wire core_csr__GEN_15 = core_csr_csr_wen & core_csr_decoded_171 &~ core_csr_reg_pmp_1_cfg_l ; 
    wire core_csr__GEN_16 = core_csr_csr_wen & core_csr_decoded_171 &~ core_csr_reg_pmp_2_cfg_l ; 
    wire core_csr__GEN_17 = core_csr_csr_wen & core_csr_decoded_171 &~ core_csr_reg_pmp_3_cfg_l ; 
    wire core_csr__GEN_18 = core_csr_csr_wen & core_csr_decoded_172 &~ core_csr_reg_pmp_4_cfg_l ; 
    wire core_csr__GEN_19 = core_csr_csr_wen & core_csr_decoded_172 &~ core_csr_reg_pmp_5_cfg_l ; 
    wire core_csr__GEN_20 = core_csr_csr_wen & core_csr_decoded_172 &~ core_csr_reg_pmp_6_cfg_l ; 
    wire core_csr__GEN_21 = core_csr_reg_pmp_7_cfg_l &~( core_csr_reg_pmp_7_cfg_a [1])& core_csr_reg_pmp_7_cfg_a [0]; 
    wire core_csr__GEN_22 = core_csr_csr_wen & core_csr_decoded_172 &~ core_csr_reg_pmp_7_cfg_l ; 
  always @( posedge  core_csr_clock )
         begin 
             if ( core_csr_reset )
                 begin  
                     core_csr_reg_mstatus_v  <=1'h0; 
                     core_csr_reg_mstatus_mpv  <=1'h0; 
                     core_csr_reg_mstatus_gva  <=1'h0; 
                     core_csr_reg_mstatus_mpp  <=2'h3; 
                     core_csr_reg_mstatus_mpie  <=1'h0; 
                     core_csr_reg_mstatus_mie  <=1'h0; 
                     core_csr_reg_dcsr_ebreakm  <=1'h0; 
                     core_csr_reg_dcsr_cause  <=3'h0; 
                     core_csr_reg_dcsr_v  <=1'h0; 
                     core_csr_reg_dcsr_step  <=1'h0; 
                     core_csr_reg_debug  <=1'h0; 
                     core_csr_reg_bp_0_control_dmode  <=1'h0; 
                     core_csr_reg_bp_0_control_action  <=1'h0; 
                     core_csr_reg_bp_0_control_x  <=1'h0; 
                     core_csr_reg_bp_0_control_w  <=1'h0; 
                     core_csr_reg_bp_0_control_r  <=1'h0; 
                     core_csr_reg_pmp_0_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_0_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_1_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_1_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_2_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_2_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_3_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_3_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_4_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_4_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_5_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_5_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_6_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_6_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_7_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_7_cfg_a  <=2'h0; 
                     core_csr_reg_mcause  <=32'h0; 
                     core_csr_reg_mtvec  <=32'h0; 
                     core_csr_reg_mcountinhibit  <=3'h0; 
                     core_csr_small_0  <=6'h0; 
                     core_csr_large_0  <=58'h0; 
                     core_csr_reg_misa  <=32'h40801105; 
                     core_csr_reg_custom_0  <=32'h8; 
                     core_csr_io_status_cease_r  <=1'h0;
                 end 
              else 
                 begin  
                     core_csr_reg_mstatus_v  <=~ core_csr_insn_ret &(~ core_csr_exception | core_csr_trapToDebug & core_csr_reg_debug )& core_csr_reg_mstatus_v ; 
                     core_csr_reg_mstatus_mpv  <= core_csr__GEN_9 &( core_csr__GEN_11  ?  core_csr_reg_mstatus_mpv : core_csr_reg_mstatus_v );
                     if ( core_csr__GEN_11 )
                         begin 
                         end 
                      else  
                         core_csr_reg_mstatus_gva  <= core_csr_io_gva ;
                     if ( core_csr__GEN_9 & core_csr__GEN_11 )
                         begin 
                         end 
                      else  
                         core_csr_reg_mstatus_mpp  <=2'h3;
                     if ( core_csr_csr_wen & core_csr_decoded_5 )
                         begin  
                             core_csr_reg_mstatus_mpie  <= core_csr_new_mstatus_mpie ; 
                             core_csr_reg_mstatus_mie  <= core_csr_new_mstatus_mie ;
                         end 
                      else 
                         begin  
                             core_csr_reg_mstatus_mpie  <= core_csr_insn_ret &~ core_csr__GEN_6 |( core_csr__GEN_11  ?  core_csr_reg_mstatus_mpie : core_csr_reg_mstatus_mie );
                             if ( core_csr__GEN_9 ) 
                                 core_csr_reg_mstatus_mie  <= core_csr__GEN_11 & core_csr_reg_mstatus_mie ;
                              else  
                                 core_csr_reg_mstatus_mie  <= core_csr_reg_mstatus_mpie ;
                         end 
                     if ( core_csr_csr_wen & core_csr_decoded_14 )
                         begin  
                             core_csr_reg_dcsr_ebreakm  <= core_csr_new_dcsr_ebreakm ; 
                             core_csr_reg_dcsr_step  <= core_csr_new_dcsr_step ;
                         end 
                     if ( core_csr__GEN_10 )
                         begin  
                             core_csr_reg_dcsr_cause  <= core_csr_reg_singleStepped  ? 3'h4:{1'h0, core_csr_causeIsDebugInt  ? 2'h3: core_csr_causeIsDebugTrigger  ? 2'h2:2'h1}; 
                             core_csr_reg_dcsr_v  <= core_csr_reg_mstatus_v ;
                         end  
                     core_csr_reg_debug  <=~( core_csr_insn_ret & core_csr__GEN_6 )&( core_csr__GEN_10 | core_csr_reg_debug );
                     if ( core_csr__GEN_13 )
                         begin  
                             core_csr_reg_bp_0_control_dmode  <= core_csr_dMode ; 
                             core_csr_reg_bp_0_control_action  <= core_csr_dMode & core_csr_newBPC_action ; 
                             core_csr_reg_bp_0_control_x  <= core_csr_wdata [2]; 
                             core_csr_reg_bp_0_control_w  <= core_csr_wdata [1]; 
                             core_csr_reg_bp_0_control_r  <= core_csr_wdata [0];
                         end 
                     if ( core_csr__GEN_14 )
                         begin  
                             core_csr_reg_pmp_0_cfg_l  <= core_csr_newCfg_l ; 
                             core_csr_reg_pmp_0_cfg_a  <= core_csr_newCfg_a ;
                         end 
                     if ( core_csr__GEN_15 )
                         begin  
                             core_csr_reg_pmp_1_cfg_l  <= core_csr_newCfg_1_l ; 
                             core_csr_reg_pmp_1_cfg_a  <= core_csr_newCfg_1_a ;
                         end 
                     if ( core_csr__GEN_16 )
                         begin  
                             core_csr_reg_pmp_2_cfg_l  <= core_csr_newCfg_2_l ; 
                             core_csr_reg_pmp_2_cfg_a  <= core_csr_newCfg_2_a ;
                         end 
                     if ( core_csr__GEN_17 )
                         begin  
                             core_csr_reg_pmp_3_cfg_l  <= core_csr_newCfg_3_l ; 
                             core_csr_reg_pmp_3_cfg_a  <= core_csr_newCfg_3_a ;
                         end 
                     if ( core_csr__GEN_18 )
                         begin  
                             core_csr_reg_pmp_4_cfg_l  <= core_csr_newCfg_4_l ; 
                             core_csr_reg_pmp_4_cfg_a  <= core_csr_newCfg_4_a ;
                         end 
                     if ( core_csr__GEN_19 )
                         begin  
                             core_csr_reg_pmp_5_cfg_l  <= core_csr_newCfg_5_l ; 
                             core_csr_reg_pmp_5_cfg_a  <= core_csr_newCfg_5_a ;
                         end 
                     if ( core_csr__GEN_20 )
                         begin  
                             core_csr_reg_pmp_6_cfg_l  <= core_csr_newCfg_6_l ; 
                             core_csr_reg_pmp_6_cfg_a  <= core_csr_newCfg_6_a ;
                         end 
                     if ( core_csr__GEN_22 )
                         begin  
                             core_csr_reg_pmp_7_cfg_l  <= core_csr_newCfg_7_l ; 
                             core_csr_reg_pmp_7_cfg_a  <= core_csr_newCfg_7_a ;
                         end 
                     if ( core_csr_csr_wen & core_csr_decoded_12 ) 
                         core_csr_reg_mcause  <= core_csr_wdata &32'h8000000F;
                      else 
                         if ( core_csr__GEN_11 )
                             begin 
                             end 
                          else  
                             core_csr_reg_mcause  <= core_csr_cause ;
                     if ( core_csr_csr_wen & core_csr_decoded_6 ) 
                         core_csr_reg_mtvec  <= core_csr_wdata ;
                     if ( core_csr_csr_wen & core_csr_decoded_17 ) 
                         core_csr_reg_mcountinhibit  <= core_csr_wdata [2:0]&3'h5;
                     if ( core_csr_csr_wen )
                         begin 
                             if ( core_csr_decoded_168 )
                                 begin  
                                     core_csr_small_0  <= core_csr_value [5:0]; 
                                     core_csr_large_0  <={ core_csr_wdata , core_csr_value [31:6]};
                                 end 
                              else 
                                 if ( core_csr_decoded_19 )
                                     begin  
                                         core_csr_small_0  <= core_csr_wdata [5:0]; 
                                         core_csr_large_0  <={ core_csr_value [63:32], core_csr_wdata [31:6]};
                                     end 
                                  else 
                                     begin 
                                         if ( core_csr_x3 )
                                             begin 
                                             end 
                                          else  
                                             core_csr_small_0  <= core_csr_nextSmall [5:0];
                                         if ( core_csr__large_T_2 ) 
                                             core_csr_large_0  <= core_csr__large_r_T ;
                                     end 
                         end 
                      else 
                         begin 
                             if ( core_csr_x3 )
                                 begin 
                                 end 
                              else  
                                 core_csr_small_0  <= core_csr_nextSmall [5:0];
                             if ( core_csr__large_T_2 ) 
                                 core_csr_large_0  <= core_csr__large_r_T ;
                         end 
                     if ( core_csr_csr_wen & core_csr_decoded_4 &(~( core_csr_io_pc [1])| core_csr_wdata [2])) 
                         core_csr_reg_misa  <=~{ core_csr__reg_misa_T [31:4], core_csr__reg_misa_T [3:0]|{~ core_csr_f ,3'h0}}&32'h1005| core_csr_reg_misa &32'hFFFFEFFA;
                     if ( core_csr_csr_wen & core_csr_decoded_191 ) 
                         core_csr_reg_custom_0  <= core_csr_wdata &32'h8| core_csr_reg_custom_0 &32'hFFFFFFF7; 
                     core_csr_io_status_cease_r  <= core_csr_insn_cease | core_csr_io_status_cease_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_15 ) 
                 core_csr_reg_dpc  <={ core_csr_wdata [31:1],1'h0};
              else 
                 if ( core_csr__GEN_10 ) 
                     core_csr_reg_dpc  <= core_csr_epc ;
             if ( core_csr_csr_wen & core_csr_decoded_16 ) 
                 core_csr_reg_dscratch0  <= core_csr_wdata ; 
             core_csr_reg_singleStepped  <= core_csr__io_singleStep_output &( core_csr_io_retire | core_csr_exception | core_csr_reg_singleStepped );
             if ( core_csr__GEN_13 ) 
                 core_csr_reg_bp_0_control_tmatch  <= core_csr_wdata [8:7];
             if ( core_csr_csr_wen & core_csr__GEN_12 & core_csr_decoded_2 ) 
                 core_csr_reg_bp_0_address  <= core_csr_wdata ;
             if ( core_csr__GEN_14 )
                 begin  
                     core_csr_reg_pmp_0_cfg_x  <= core_csr_newCfg_x ; 
                     core_csr_reg_pmp_0_cfg_w  <= core_csr_newCfg_w & core_csr_newCfg_r ; 
                     core_csr_reg_pmp_0_cfg_r  <= core_csr_newCfg_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_175 &~( core_csr_reg_pmp_0_cfg_l | core_csr_reg_pmp_1_cfg_l &~( core_csr_reg_pmp_1_cfg_a [1])& core_csr_reg_pmp_1_cfg_a [0])) 
                 core_csr_reg_pmp_0_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_15 )
                 begin  
                     core_csr_reg_pmp_1_cfg_x  <= core_csr_newCfg_1_x ; 
                     core_csr_reg_pmp_1_cfg_w  <= core_csr_newCfg_1_w & core_csr_newCfg_1_r ; 
                     core_csr_reg_pmp_1_cfg_r  <= core_csr_newCfg_1_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_176 &~( core_csr_reg_pmp_1_cfg_l | core_csr_reg_pmp_2_cfg_l &~( core_csr_reg_pmp_2_cfg_a [1])& core_csr_reg_pmp_2_cfg_a [0])) 
                 core_csr_reg_pmp_1_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_16 )
                 begin  
                     core_csr_reg_pmp_2_cfg_x  <= core_csr_newCfg_2_x ; 
                     core_csr_reg_pmp_2_cfg_w  <= core_csr_newCfg_2_w & core_csr_newCfg_2_r ; 
                     core_csr_reg_pmp_2_cfg_r  <= core_csr_newCfg_2_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_177 &~( core_csr_reg_pmp_2_cfg_l | core_csr_reg_pmp_3_cfg_l &~( core_csr_reg_pmp_3_cfg_a [1])& core_csr_reg_pmp_3_cfg_a [0])) 
                 core_csr_reg_pmp_2_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_17 )
                 begin  
                     core_csr_reg_pmp_3_cfg_x  <= core_csr_newCfg_3_x ; 
                     core_csr_reg_pmp_3_cfg_w  <= core_csr_newCfg_3_w & core_csr_newCfg_3_r ; 
                     core_csr_reg_pmp_3_cfg_r  <= core_csr_newCfg_3_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_178 &~( core_csr_reg_pmp_3_cfg_l | core_csr_reg_pmp_4_cfg_l &~( core_csr_reg_pmp_4_cfg_a [1])& core_csr_reg_pmp_4_cfg_a [0])) 
                 core_csr_reg_pmp_3_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_18 )
                 begin  
                     core_csr_reg_pmp_4_cfg_x  <= core_csr_newCfg_4_x ; 
                     core_csr_reg_pmp_4_cfg_w  <= core_csr_newCfg_4_w & core_csr_newCfg_4_r ; 
                     core_csr_reg_pmp_4_cfg_r  <= core_csr_newCfg_4_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_179 &~( core_csr_reg_pmp_4_cfg_l | core_csr_reg_pmp_5_cfg_l &~( core_csr_reg_pmp_5_cfg_a [1])& core_csr_reg_pmp_5_cfg_a [0])) 
                 core_csr_reg_pmp_4_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_19 )
                 begin  
                     core_csr_reg_pmp_5_cfg_x  <= core_csr_newCfg_5_x ; 
                     core_csr_reg_pmp_5_cfg_w  <= core_csr_newCfg_5_w & core_csr_newCfg_5_r ; 
                     core_csr_reg_pmp_5_cfg_r  <= core_csr_newCfg_5_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_180 &~( core_csr_reg_pmp_5_cfg_l | core_csr_reg_pmp_6_cfg_l &~( core_csr_reg_pmp_6_cfg_a [1])& core_csr_reg_pmp_6_cfg_a [0])) 
                 core_csr_reg_pmp_5_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_20 )
                 begin  
                     core_csr_reg_pmp_6_cfg_x  <= core_csr_newCfg_6_x ; 
                     core_csr_reg_pmp_6_cfg_w  <= core_csr_newCfg_6_w & core_csr_newCfg_6_r ; 
                     core_csr_reg_pmp_6_cfg_r  <= core_csr_newCfg_6_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_181 &~( core_csr_reg_pmp_6_cfg_l | core_csr__GEN_21 )) 
                 core_csr_reg_pmp_6_addr  <= core_csr_wdata [29:0];
             if ( core_csr__GEN_22 )
                 begin  
                     core_csr_reg_pmp_7_cfg_x  <= core_csr_newCfg_7_x ; 
                     core_csr_reg_pmp_7_cfg_w  <= core_csr_newCfg_7_w & core_csr_newCfg_7_r ; 
                     core_csr_reg_pmp_7_cfg_r  <= core_csr_newCfg_7_r ;
                 end 
             if ( core_csr_csr_wen & core_csr_decoded_182 &~( core_csr_reg_pmp_7_cfg_l | core_csr__GEN_21 )) 
                 core_csr_reg_pmp_7_addr  <= core_csr_wdata [29:0];
             if ( core_csr_csr_wen & core_csr_decoded_8 ) 
                 core_csr_reg_mie  <={20'h0, core_csr_wdata [11:3]&9'h111,3'h0};
             if ( core_csr_csr_wen & core_csr_decoded_10 ) 
                 core_csr_reg_mepc  <={ core_csr_wdata [31:1],1'h0};
              else 
                 if ( core_csr__GEN_11 )
                     begin 
                     end 
                  else  
                     core_csr_reg_mepc  <= core_csr_epc ;
             if ( core_csr_csr_wen & core_csr_decoded_11 ) 
                 core_csr_reg_mtval  <= core_csr_wdata ;
              else 
                 if ( core_csr__GEN_11 )
                     begin 
                     end 
                  else  
                     core_csr_reg_mtval  <= core_csr_tval ;
             if ( core_csr__GEN_11 )
                 begin 
                 end 
              else  
                 core_csr_reg_mtval2  <= core_csr_io_htval ;
             if ( core_csr_csr_wen & core_csr_decoded_9 ) 
                 core_csr_reg_mscratch  <= core_csr_wdata ;
         end
    wire core_csr__large_T_5 = core_csr_nextSmall_1 [6]&~ core_csr_x11 ; 
    wire[57:0] core_csr__large_r_T_2 = core_csr_large_1 +58'h1; 
  always @( posedge  core_csr_io_ungated_clock )
         begin 
             if ( core_csr_reset )
                 begin  
                     core_csr_reg_wfi  <=1'h0; 
                     core_csr_small_1  <=6'h0; 
                     core_csr_large_1  <=58'h0;
                 end 
              else 
                 begin  
                     core_csr_reg_wfi  <=~((| core_csr_pending_interrupts )| core_csr_io_interrupts_debug | core_csr_exception )&( core_csr_insn_wfi &~ core_csr__io_singleStep_output &~ core_csr_reg_debug | core_csr_reg_wfi );
                     if ( core_csr_csr_wen )
                         begin 
                             if ( core_csr_decoded_167 )
                                 begin  
                                     core_csr_small_1  <= core_csr_value_1 [5:0]; 
                                     core_csr_large_1  <={ core_csr_wdata , core_csr_value_1 [31:6]};
                                 end 
                              else 
                                 if ( core_csr_decoded_18 )
                                     begin  
                                         core_csr_small_1  <= core_csr_wdata [5:0]; 
                                         core_csr_large_1  <={ core_csr_value_1 [63:32], core_csr_wdata [31:6]};
                                     end 
                                  else 
                                     begin 
                                         if ( core_csr_x11 )
                                             begin 
                                             end 
                                          else  
                                             core_csr_small_1  <= core_csr_nextSmall_1 [5:0];
                                         if ( core_csr__large_T_5 ) 
                                             core_csr_large_1  <= core_csr__large_r_T_2 ;
                                     end 
                         end 
                      else 
                         begin 
                             if ( core_csr_x11 )
                                 begin 
                                 end 
                              else  
                                 core_csr_small_1  <= core_csr_nextSmall_1 [5:0];
                             if ( core_csr__large_T_5 ) 
                                 core_csr_large_1  <= core_csr__large_r_T_2 ;
                         end 
                 end 
         end
  assign  core_csr_io_rw_rdata = core_csr__io_rw_rdata_output ; 
  assign  core_csr_io_decode_0_read_illegal =~ core_csr_csr_addr_legal |~ core_csr_csr_exists | core_csr_io_decode_0_read_illegal_plaOutput &~ core_csr_reg_debug ; 
  assign  core_csr_io_decode_0_write_illegal =&( core_csr_addr_1 [11:10]); 
  assign  core_csr_io_decode_0_write_flush =~( core_csr_io_decode_0_write_flush_addr_m >12'h33F& core_csr_io_decode_0_write_flush_addr_m <12'h344); 
  assign  core_csr_io_decode_0_system_illegal =~ core_csr_csr_addr_legal &~ core_csr_is_hlsv | core_csr_is_ret & core_csr_addr_1 [10]& core_csr_addr_1 [7]&~ core_csr_reg_debug ; 
  assign  core_csr_io_decode_0_virtual_access_illegal = core_csr_reg_mstatus_v & core_csr_csr_exists &( core_csr_addr_1 [9:8]==2'h2| core_csr_is_counter & core_csr__io_decode_0_virtual_access_illegal_T_3 [0]&~( core_csr__io_decode_0_virtual_access_illegal_T_6 [0])); 
  assign  core_csr_io_decode_0_virtual_system_illegal = core_csr_reg_mstatus_v &( core_csr_is_hfence_vvma | core_csr_is_hfence_gvma | core_csr_is_hlsv ); 
  assign  core_csr_io_csr_stall = core_csr__io_csr_stall_output ; 
  assign  core_csr_io_eret = core_csr__exception_T | core_csr_insn_ret ; 
  assign  core_csr_io_singleStep = core_csr__io_singleStep_output ; 
  assign  core_csr_io_status_debug = core_csr_reg_debug ; 
  assign  core_csr_io_status_wfi = core_csr_reg_wfi ; 
  assign  core_csr_io_status_isa = core_csr_reg_misa ; 
  assign  core_csr_io_status_dv = core_csr_reg_mstatus_v ; 
  assign  core_csr_io_status_v = core_csr_reg_mstatus_v ; 
  assign  core_csr_io_evec = core_csr_insn_ret  ? ( core_csr__GEN_6  ? ~{ core_csr__io_evec_T_10 [31:2], core_csr__io_evec_T_10 [1:0]|{~( core_csr_reg_misa [2]),1'h1}}:~{ core_csr__io_evec_T_20 [31:2], core_csr__io_evec_T_20 [1:0]|{~( core_csr_reg_misa [2]),1'h1}}): core_csr_tvec ; 
  assign  core_csr_io_time = core_csr_value_1 [31:0]; 
  assign  core_csr_io_interrupt =( core_csr_anyInterrupt &~ core_csr__io_singleStep_output | core_csr_reg_singleStepped )&~( core_csr_reg_debug | core_csr_io_status_cease_r ); 
  assign  core_csr_io_interrupt_cause = core_csr_interruptCause ; 
  assign  core_csr_io_bp_0_control_action = core_csr_reg_bp_0_control_action ; 
  assign  core_csr_io_bp_0_control_tmatch = core_csr_reg_bp_0_control_tmatch ; 
  assign  core_csr_io_bp_0_control_x = core_csr_reg_bp_0_control_x ; 
  assign  core_csr_io_bp_0_control_w = core_csr_reg_bp_0_control_w ; 
  assign  core_csr_io_bp_0_control_r = core_csr_reg_bp_0_control_r ; 
  assign  core_csr_io_bp_0_address = core_csr_reg_bp_0_address ; 
  assign  core_csr_io_pmp_0_cfg_l = core_csr_pmp_cfg_l ; 
  assign  core_csr_io_pmp_0_cfg_a = core_csr_pmp_cfg_a ; 
  assign  core_csr_io_pmp_0_cfg_x = core_csr_pmp_cfg_x ; 
  assign  core_csr_io_pmp_0_cfg_w = core_csr_pmp_cfg_w ; 
  assign  core_csr_io_pmp_0_cfg_r = core_csr_pmp_cfg_r ; 
  assign  core_csr_io_pmp_0_addr = core_csr_pmp_addr ; 
  assign  core_csr_io_pmp_0_mask = core_csr_pmp_mask ; 
  assign  core_csr_io_pmp_1_cfg_l = core_csr_pmp_1_cfg_l ; 
  assign  core_csr_io_pmp_1_cfg_a = core_csr_pmp_1_cfg_a ; 
  assign  core_csr_io_pmp_1_cfg_x = core_csr_pmp_1_cfg_x ; 
  assign  core_csr_io_pmp_1_cfg_w = core_csr_pmp_1_cfg_w ; 
  assign  core_csr_io_pmp_1_cfg_r = core_csr_pmp_1_cfg_r ; 
  assign  core_csr_io_pmp_1_addr = core_csr_pmp_1_addr ; 
  assign  core_csr_io_pmp_1_mask = core_csr_pmp_1_mask ; 
  assign  core_csr_io_pmp_2_cfg_l = core_csr_pmp_2_cfg_l ; 
  assign  core_csr_io_pmp_2_cfg_a = core_csr_pmp_2_cfg_a ; 
  assign  core_csr_io_pmp_2_cfg_x = core_csr_pmp_2_cfg_x ; 
  assign  core_csr_io_pmp_2_cfg_w = core_csr_pmp_2_cfg_w ; 
  assign  core_csr_io_pmp_2_cfg_r = core_csr_pmp_2_cfg_r ; 
  assign  core_csr_io_pmp_2_addr = core_csr_pmp_2_addr ; 
  assign  core_csr_io_pmp_2_mask = core_csr_pmp_2_mask ; 
  assign  core_csr_io_pmp_3_cfg_l = core_csr_pmp_3_cfg_l ; 
  assign  core_csr_io_pmp_3_cfg_a = core_csr_pmp_3_cfg_a ; 
  assign  core_csr_io_pmp_3_cfg_x = core_csr_pmp_3_cfg_x ; 
  assign  core_csr_io_pmp_3_cfg_w = core_csr_pmp_3_cfg_w ; 
  assign  core_csr_io_pmp_3_cfg_r = core_csr_pmp_3_cfg_r ; 
  assign  core_csr_io_pmp_3_addr = core_csr_pmp_3_addr ; 
  assign  core_csr_io_pmp_3_mask = core_csr_pmp_3_mask ; 
  assign  core_csr_io_pmp_4_cfg_l = core_csr_pmp_4_cfg_l ; 
  assign  core_csr_io_pmp_4_cfg_a = core_csr_pmp_4_cfg_a ; 
  assign  core_csr_io_pmp_4_cfg_x = core_csr_pmp_4_cfg_x ; 
  assign  core_csr_io_pmp_4_cfg_w = core_csr_pmp_4_cfg_w ; 
  assign  core_csr_io_pmp_4_cfg_r = core_csr_pmp_4_cfg_r ; 
  assign  core_csr_io_pmp_4_addr = core_csr_pmp_4_addr ; 
  assign  core_csr_io_pmp_4_mask = core_csr_pmp_4_mask ; 
  assign  core_csr_io_pmp_5_cfg_l = core_csr_pmp_5_cfg_l ; 
  assign  core_csr_io_pmp_5_cfg_a = core_csr_pmp_5_cfg_a ; 
  assign  core_csr_io_pmp_5_cfg_x = core_csr_pmp_5_cfg_x ; 
  assign  core_csr_io_pmp_5_cfg_w = core_csr_pmp_5_cfg_w ; 
  assign  core_csr_io_pmp_5_cfg_r = core_csr_pmp_5_cfg_r ; 
  assign  core_csr_io_pmp_5_addr = core_csr_pmp_5_addr ; 
  assign  core_csr_io_pmp_5_mask = core_csr_pmp_5_mask ; 
  assign  core_csr_io_pmp_6_cfg_l = core_csr_pmp_6_cfg_l ; 
  assign  core_csr_io_pmp_6_cfg_a = core_csr_pmp_6_cfg_a ; 
  assign  core_csr_io_pmp_6_cfg_x = core_csr_pmp_6_cfg_x ; 
  assign  core_csr_io_pmp_6_cfg_w = core_csr_pmp_6_cfg_w ; 
  assign  core_csr_io_pmp_6_cfg_r = core_csr_pmp_6_cfg_r ; 
  assign  core_csr_io_pmp_6_addr = core_csr_pmp_6_addr ; 
  assign  core_csr_io_pmp_6_mask = core_csr_pmp_6_mask ; 
  assign  core_csr_io_pmp_7_cfg_l = core_csr_pmp_7_cfg_l ; 
  assign  core_csr_io_pmp_7_cfg_a = core_csr_pmp_7_cfg_a ; 
  assign  core_csr_io_pmp_7_cfg_x = core_csr_pmp_7_cfg_x ; 
  assign  core_csr_io_pmp_7_cfg_w = core_csr_pmp_7_cfg_w ; 
  assign  core_csr_io_pmp_7_cfg_r = core_csr_pmp_7_cfg_r ; 
  assign  core_csr_io_pmp_7_addr = core_csr_pmp_7_addr ; 
  assign  core_csr_io_pmp_7_mask = core_csr_pmp_7_mask ; 
  assign  core_csr_io_inhibit_cycle = core_csr_x11 ; 
  assign  core_csr_io_trace_0_valid = core_csr_io_retire | core_csr_exception ; 
  assign  core_csr_io_trace_0_iaddr = core_csr_io_pc ; 
  assign  core_csr_io_trace_0_insn = core_csr_io_inst_0 ; 
  assign  core_csr_io_trace_0_priv ={ core_csr_reg_debug ,2'h3}; 
  assign  core_csr_io_trace_0_exception = core_csr_exception ; 
  assign  core_csr_io_trace_0_interrupt = core_csr_cause [31]; 
  assign  core_csr_io_trace_0_cause = core_csr_cause ; 
  assign  core_csr_io_trace_0_tval = core_csr_io_tval ; 
  assign  core_csr_io_customCSRs_0_value = core_csr_reg_custom_0 ;
    assign core_csr_clock = core_clock;
    assign core_csr_reset = core_reset;
    assign core_csr_io_ungated_clock = core_clock;
    assign core_csr_io_interrupts_debug = core_io_interrupts_debug;
    assign core_csr_io_interrupts_mtip = core_io_interrupts_mtip;
    assign core_csr_io_interrupts_msip = core_io_interrupts_msip;
    assign core_csr_io_interrupts_meip = core_io_interrupts_meip;
    assign core_csr_io_hartid = core_io_hartid;
    assign core_csr_io_rw_addr = core_wb_reg_inst[31:20];
    assign core_csr_io_rw_cmd = core_wb_ctrl_csr&{core_wb_reg_valid,2'h3};
    assign core__csr_io_rw_rdata = core_csr_io_rw_rdata;
    assign core_csr_io_rw_wdata = core_wb_reg_wdata;
    assign core_csr_io_decode_0_inst = core__ibuf_io_inst_0_bits_inst_bits;
    assign core__csr_io_decode_0_read_illegal = core_csr_io_decode_0_read_illegal;
    assign core__csr_io_decode_0_write_illegal = core_csr_io_decode_0_write_illegal;
    assign core__csr_io_decode_0_write_flush = core_csr_io_decode_0_write_flush;
    assign core__csr_io_decode_0_system_illegal = core_csr_io_decode_0_system_illegal;
    assign core__csr_io_decode_0_virtual_access_illegal = core_csr_io_decode_0_virtual_access_illegal;
    assign core__csr_io_decode_0_virtual_system_illegal = core_csr_io_decode_0_virtual_system_illegal;
    assign core__csr_io_csr_stall = core_csr_io_csr_stall;
    assign core__csr_io_eret = core_csr_io_eret;
    assign core__csr_io_singleStep = core_csr_io_singleStep;
    assign core__csr_io_status_debug = core_csr_io_status_debug;
    assign core_io_wfi = core_csr_io_status_wfi;
    assign core__csr_io_status_isa = core_csr_io_status_isa;
    assign core__csr_io_status_dv = core_csr_io_status_dv;
    assign core__csr_io_status_v = core_csr_io_status_v;
    assign core__csr_io_evec = core_csr_io_evec;
    assign core_csr_io_exception = core_wb_xcpt;
    assign core_csr_io_retire = core_wb_valid;
    assign core_csr_io_cause = core_wb_cause;
    assign core_csr_io_pc = core_wb_reg_pc;
    assign core_csr_io_tval = core_tval_valid ? core_wb_reg_wdata:32'h0;
    assign core_csr_io_htval = core_csr_io_htval_htval_imem;
    assign core_csr_io_gva = core_wb_xcpt&(core_tval_any_addr&core__csr_io_status_v|core_tval_dmem_addr&core_wb_reg_hls_or_dv);
    assign core__csr_io_time = core_csr_io_time;
    assign core__csr_io_interrupt = core_csr_io_interrupt;
    assign core__csr_io_interrupt_cause = core_csr_io_interrupt_cause;
    assign core__csr_io_bp_0_control_action = core_csr_io_bp_0_control_action;
    assign core__csr_io_bp_0_control_tmatch = core_csr_io_bp_0_control_tmatch;
    assign core__csr_io_bp_0_control_x = core_csr_io_bp_0_control_x;
    assign core__csr_io_bp_0_control_w = core_csr_io_bp_0_control_w;
    assign core__csr_io_bp_0_control_r = core_csr_io_bp_0_control_r;
    assign core__csr_io_bp_0_address = core_csr_io_bp_0_address;
    assign core_io_ptw_pmp_0_cfg_l = core_csr_io_pmp_0_cfg_l;
    assign core_io_ptw_pmp_0_cfg_a = core_csr_io_pmp_0_cfg_a;
    assign core_io_ptw_pmp_0_cfg_x = core_csr_io_pmp_0_cfg_x;
    assign core_io_ptw_pmp_0_cfg_w = core_csr_io_pmp_0_cfg_w;
    assign core_io_ptw_pmp_0_cfg_r = core_csr_io_pmp_0_cfg_r;
    assign core_io_ptw_pmp_0_addr = core_csr_io_pmp_0_addr;
    assign core_io_ptw_pmp_0_mask = core_csr_io_pmp_0_mask;
    assign core_io_ptw_pmp_1_cfg_l = core_csr_io_pmp_1_cfg_l;
    assign core_io_ptw_pmp_1_cfg_a = core_csr_io_pmp_1_cfg_a;
    assign core_io_ptw_pmp_1_cfg_x = core_csr_io_pmp_1_cfg_x;
    assign core_io_ptw_pmp_1_cfg_w = core_csr_io_pmp_1_cfg_w;
    assign core_io_ptw_pmp_1_cfg_r = core_csr_io_pmp_1_cfg_r;
    assign core_io_ptw_pmp_1_addr = core_csr_io_pmp_1_addr;
    assign core_io_ptw_pmp_1_mask = core_csr_io_pmp_1_mask;
    assign core_io_ptw_pmp_2_cfg_l = core_csr_io_pmp_2_cfg_l;
    assign core_io_ptw_pmp_2_cfg_a = core_csr_io_pmp_2_cfg_a;
    assign core_io_ptw_pmp_2_cfg_x = core_csr_io_pmp_2_cfg_x;
    assign core_io_ptw_pmp_2_cfg_w = core_csr_io_pmp_2_cfg_w;
    assign core_io_ptw_pmp_2_cfg_r = core_csr_io_pmp_2_cfg_r;
    assign core_io_ptw_pmp_2_addr = core_csr_io_pmp_2_addr;
    assign core_io_ptw_pmp_2_mask = core_csr_io_pmp_2_mask;
    assign core_io_ptw_pmp_3_cfg_l = core_csr_io_pmp_3_cfg_l;
    assign core_io_ptw_pmp_3_cfg_a = core_csr_io_pmp_3_cfg_a;
    assign core_io_ptw_pmp_3_cfg_x = core_csr_io_pmp_3_cfg_x;
    assign core_io_ptw_pmp_3_cfg_w = core_csr_io_pmp_3_cfg_w;
    assign core_io_ptw_pmp_3_cfg_r = core_csr_io_pmp_3_cfg_r;
    assign core_io_ptw_pmp_3_addr = core_csr_io_pmp_3_addr;
    assign core_io_ptw_pmp_3_mask = core_csr_io_pmp_3_mask;
    assign core_io_ptw_pmp_4_cfg_l = core_csr_io_pmp_4_cfg_l;
    assign core_io_ptw_pmp_4_cfg_a = core_csr_io_pmp_4_cfg_a;
    assign core_io_ptw_pmp_4_cfg_x = core_csr_io_pmp_4_cfg_x;
    assign core_io_ptw_pmp_4_cfg_w = core_csr_io_pmp_4_cfg_w;
    assign core_io_ptw_pmp_4_cfg_r = core_csr_io_pmp_4_cfg_r;
    assign core_io_ptw_pmp_4_addr = core_csr_io_pmp_4_addr;
    assign core_io_ptw_pmp_4_mask = core_csr_io_pmp_4_mask;
    assign core_io_ptw_pmp_5_cfg_l = core_csr_io_pmp_5_cfg_l;
    assign core_io_ptw_pmp_5_cfg_a = core_csr_io_pmp_5_cfg_a;
    assign core_io_ptw_pmp_5_cfg_x = core_csr_io_pmp_5_cfg_x;
    assign core_io_ptw_pmp_5_cfg_w = core_csr_io_pmp_5_cfg_w;
    assign core_io_ptw_pmp_5_cfg_r = core_csr_io_pmp_5_cfg_r;
    assign core_io_ptw_pmp_5_addr = core_csr_io_pmp_5_addr;
    assign core_io_ptw_pmp_5_mask = core_csr_io_pmp_5_mask;
    assign core_io_ptw_pmp_6_cfg_l = core_csr_io_pmp_6_cfg_l;
    assign core_io_ptw_pmp_6_cfg_a = core_csr_io_pmp_6_cfg_a;
    assign core_io_ptw_pmp_6_cfg_x = core_csr_io_pmp_6_cfg_x;
    assign core_io_ptw_pmp_6_cfg_w = core_csr_io_pmp_6_cfg_w;
    assign core_io_ptw_pmp_6_cfg_r = core_csr_io_pmp_6_cfg_r;
    assign core_io_ptw_pmp_6_addr = core_csr_io_pmp_6_addr;
    assign core_io_ptw_pmp_6_mask = core_csr_io_pmp_6_mask;
    assign core_io_ptw_pmp_7_cfg_l = core_csr_io_pmp_7_cfg_l;
    assign core_io_ptw_pmp_7_cfg_a = core_csr_io_pmp_7_cfg_a;
    assign core_io_ptw_pmp_7_cfg_x = core_csr_io_pmp_7_cfg_x;
    assign core_io_ptw_pmp_7_cfg_w = core_csr_io_pmp_7_cfg_w;
    assign core_io_ptw_pmp_7_cfg_r = core_csr_io_pmp_7_cfg_r;
    assign core_io_ptw_pmp_7_addr = core_csr_io_pmp_7_addr;
    assign core_io_ptw_pmp_7_mask = core_csr_io_pmp_7_mask;
    assign core__csr_io_inhibit_cycle = core_csr_io_inhibit_cycle;
    assign core_csr_io_inst_0 = {(&(core_wb_reg_raw_inst[1:0])) ? core_wb_reg_inst[31:16]:16'h0,core_wb_reg_raw_inst[15:0]};
    assign core__csr_io_trace_0_valid = core_csr_io_trace_0_valid;
    assign core__csr_io_trace_0_iaddr = core_csr_io_trace_0_iaddr;
    assign core__csr_io_trace_0_insn = core_csr_io_trace_0_insn;
    assign core__csr_io_trace_0_priv = core_csr_io_trace_0_priv;
    assign core__csr_io_trace_0_exception = core_csr_io_trace_0_exception;
    assign core_io_trace_insns_0_interrupt = core_csr_io_trace_0_interrupt;
    assign core_io_trace_insns_0_cause = core_csr_io_trace_0_cause;
    assign core_io_trace_insns_0_tval = core_csr_io_trace_0_tval;
    assign core__csr_io_customCSRs_0_value = core_csr_io_customCSRs_0_value;
     
    wire core_coreMonitorBundle_excpt ; 
  assign  core_coreMonitorBundle_excpt = core__csr_io_trace_0_exception ; 
    wire[2:0] core_coreMonitorBundle_priv_mode ; 
  assign  core_coreMonitorBundle_priv_mode = core__csr_io_trace_0_priv ; 
  assign  core_coreMonitorBundle_timer = core__csr_io_time ; 
  assign  core_coreMonitorBundle_pc = core__csr_io_trace_0_iaddr ; 
  assign  core_coreMonitorBundle_inst = core__csr_io_trace_0_insn ; 
    wire[2:0] core_xrfWriteBundle_priv_mode ; 
  assign  core_xrfWriteBundle_priv_mode = core__csr_io_trace_0_priv ; 
    wire[31:0] core_xrfWriteBundle_timer ; 
  assign  core_xrfWriteBundle_timer = core__csr_io_time ;  
    wire core_bpu_io_status_debug;
    wire core_bpu_io_bp_0_control_action;
    wire[1:0] core_bpu_io_bp_0_control_tmatch;
    wire core_bpu_io_bp_0_control_x;
    wire core_bpu_io_bp_0_control_w;
    wire core_bpu_io_bp_0_control_r;
    wire[31:0] core_bpu_io_bp_0_address;
    wire[31:0] core_bpu_io_pc;
    wire[31:0] core_bpu_io_ea;
    wire core_bpu_io_xcpt_if;
    wire core_bpu_io_xcpt_ld;
    wire core_bpu_io_xcpt_st;
    wire core_bpu_io_debug_if;
    wire core_bpu_io_debug_ld;
    wire core_bpu_io_debug_st;
    wire core_bpu_io_bpwatch_0_rvalid_0;
    wire core_bpu_io_bpwatch_0_wvalid_0;
    wire core_bpu_io_bpwatch_0_ivalid_0;

    wire[1:0] core_bpu_en_lo =2'h0; 
    wire[1:0] core_bpu_en_hi =2'h2; 
    wire core_bpu_cx =1'h1; 
    wire core_bpu_end_0 =1'h1; 
    wire core_bpu_en =~ core_bpu_io_status_debug ; 
    wire core_bpu__w_T_2 = core_bpu_io_ea >= core_bpu_io_bp_0_address ; 
    wire[31:0] core_bpu__w_T_5 =~ core_bpu_io_ea ; 
    wire core_bpu__r_T_8 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__r_T_10 = core_bpu__r_T_8 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_r_lo ={ core_bpu__r_T_8 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_r_hi ={ core_bpu__r_T_10 & core_bpu_io_bp_0_address [2], core_bpu__r_T_10 }; 
    wire[31:0] core_bpu__x_T_15 =~ core_bpu_io_bp_0_address ; 
    wire core_bpu__r_T_18 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__r_T_20 = core_bpu__r_T_18 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_r_lo_1 ={ core_bpu__r_T_18 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_r_hi_1 ={ core_bpu__r_T_20 & core_bpu_io_bp_0_address [2], core_bpu__r_T_20 }; 
    wire core_bpu_r = core_bpu_en & core_bpu_io_bp_0_control_r &( core_bpu_io_bp_0_control_tmatch [1] ?  core_bpu__w_T_2 ^ core_bpu_io_bp_0_control_tmatch [0]:{ core_bpu__w_T_5 [31:4], core_bpu__w_T_5 [3:0]|{ core_bpu_r_hi , core_bpu_r_lo }}=={ core_bpu__x_T_15 [31:4], core_bpu__x_T_15 [3:0]|{ core_bpu_r_hi_1 , core_bpu_r_lo_1 }}); 
    wire core_bpu__w_T_8 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__w_T_10 = core_bpu__w_T_8 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_w_lo ={ core_bpu__w_T_8 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_w_hi ={ core_bpu__w_T_10 & core_bpu_io_bp_0_address [2], core_bpu__w_T_10 }; 
    wire core_bpu__w_T_18 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__w_T_20 = core_bpu__w_T_18 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_w_lo_1 ={ core_bpu__w_T_18 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_w_hi_1 ={ core_bpu__w_T_20 & core_bpu_io_bp_0_address [2], core_bpu__w_T_20 }; 
    wire core_bpu_w = core_bpu_en & core_bpu_io_bp_0_control_w &( core_bpu_io_bp_0_control_tmatch [1] ?  core_bpu__w_T_2 ^ core_bpu_io_bp_0_control_tmatch [0]:{ core_bpu__w_T_5 [31:4], core_bpu__w_T_5 [3:0]|{ core_bpu_w_hi , core_bpu_w_lo }}=={ core_bpu__x_T_15 [31:4], core_bpu__x_T_15 [3:0]|{ core_bpu_w_hi_1 , core_bpu_w_lo_1 }}); 
    wire[31:0] core_bpu__x_T_5 =~ core_bpu_io_pc ; 
    wire core_bpu__x_T_8 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__x_T_10 = core_bpu__x_T_8 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_x_lo ={ core_bpu__x_T_8 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_x_hi ={ core_bpu__x_T_10 & core_bpu_io_bp_0_address [2], core_bpu__x_T_10 }; 
    wire core_bpu__x_T_18 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__x_T_20 = core_bpu__x_T_18 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_x_lo_1 ={ core_bpu__x_T_18 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_x_hi_1 ={ core_bpu__x_T_20 & core_bpu_io_bp_0_address [2], core_bpu__x_T_20 }; 
    wire core_bpu_x = core_bpu_en & core_bpu_io_bp_0_control_x &( core_bpu_io_bp_0_control_tmatch [1] ?  core_bpu_io_pc >= core_bpu_io_bp_0_address ^ core_bpu_io_bp_0_control_tmatch [0]:{ core_bpu__x_T_5 [31:4], core_bpu__x_T_5 [3:0]|{ core_bpu_x_hi , core_bpu_x_lo }}=={ core_bpu__x_T_15 [31:4], core_bpu__x_T_15 [3:0]|{ core_bpu_x_hi_1 , core_bpu_x_lo_1 }}); 
  assign  core_bpu_io_xcpt_if = core_bpu_x &~ core_bpu_io_bp_0_control_action ; 
  assign  core_bpu_io_xcpt_ld = core_bpu_r &~ core_bpu_io_bp_0_control_action ; 
  assign  core_bpu_io_xcpt_st = core_bpu_w &~ core_bpu_io_bp_0_control_action ; 
  assign  core_bpu_io_debug_if = core_bpu_x & core_bpu_io_bp_0_control_action ; 
  assign  core_bpu_io_debug_ld = core_bpu_r & core_bpu_io_bp_0_control_action ; 
  assign  core_bpu_io_debug_st = core_bpu_w & core_bpu_io_bp_0_control_action ; 
  assign  core_bpu_io_bpwatch_0_rvalid_0 = core_bpu_r ; 
  assign  core_bpu_io_bpwatch_0_wvalid_0 = core_bpu_w ; 
  assign  core_bpu_io_bpwatch_0_ivalid_0 = core_bpu_x ;
    assign core_bpu_io_status_debug = core__csr_io_status_debug;
    assign core_bpu_io_bp_0_control_action = core__csr_io_bp_0_control_action;
    assign core_bpu_io_bp_0_control_tmatch = core__csr_io_bp_0_control_tmatch;
    assign core_bpu_io_bp_0_control_x = core__csr_io_bp_0_control_x;
    assign core_bpu_io_bp_0_control_w = core__csr_io_bp_0_control_w;
    assign core_bpu_io_bp_0_control_r = core__csr_io_bp_0_control_r;
    assign core_bpu_io_bp_0_address = core__csr_io_bp_0_address;
    assign core_bpu_io_pc = core__ibuf_io_pc;
    assign core_bpu_io_ea = core_mem_reg_wdata;
    assign core__bpu_io_xcpt_if = core_bpu_io_xcpt_if;
    assign core__bpu_io_xcpt_ld = core_bpu_io_xcpt_ld;
    assign core__bpu_io_xcpt_st = core_bpu_io_xcpt_st;
    assign core__bpu_io_debug_if = core_bpu_io_debug_if;
    assign core__bpu_io_debug_ld = core_bpu_io_debug_ld;
    assign core__bpu_io_debug_st = core_bpu_io_debug_st;
    assign core__bpu_io_bpwatch_0_rvalid_0 = core_bpu_io_bpwatch_0_rvalid_0;
    assign core__bpu_io_bpwatch_0_wvalid_0 = core_bpu_io_bpwatch_0_wvalid_0;
    assign core__bpu_io_bpwatch_0_ivalid_0 = core_bpu_io_bpwatch_0_ivalid_0;
      
    wire[3:0] core_alu_io_fn;
    wire[31:0] core_alu_io_in2;
    wire[31:0] core_alu_io_in1;
    wire[31:0] core_alu_io_out;
    wire[31:0] core_alu_io_adder_out;
    wire core_alu_io_cmp_out;

    wire[31:0] core_alu_in2_inv ={32{ core_alu_io_fn [3]}}^ core_alu_io_in2 ; 
    wire[31:0] core_alu_in1_xor_in2 = core_alu_io_in1 ^ core_alu_in2_inv ; 
    wire[31:0] core_alu__io_adder_out_T_3 = core_alu_io_in1 + core_alu_in2_inv +{31'h0, core_alu_io_fn [3]}; 
    wire core_alu_slt = core_alu_io_in1 [31]== core_alu_io_in2 [31] ?  core_alu__io_adder_out_T_3 [31]: core_alu_io_fn [1] ?  core_alu_io_in2 [31]: core_alu_io_in1 [31]; 
    wire[4:0] core_alu_shamt = core_alu_io_in2 [4:0]; 
    wire core_alu__shout_T = core_alu_io_fn ==4'h5; 
    wire core_alu__shout_T_1 = core_alu_io_fn ==4'hB; 
    wire[7:0] core_alu__GEN ={{ core_alu_io_in1 [11:8], core_alu_io_in1 [15:14]}&6'h33,2'h0}|{ core_alu_io_in1 [15:12], core_alu_io_in1 [19:16]}&8'h33; 
    wire[18:0] core_alu__GEN_0 ={ core_alu_io_in1 [5:4], core_alu_io_in1 [7:6], core_alu_io_in1 [9:8], core_alu__GEN , core_alu_io_in1 [19:18], core_alu_io_in1 [21:20], core_alu_io_in1 [23]}&19'h55555; 
    wire[31:0] core_alu_shin = core_alu__shout_T | core_alu__shout_T_1  ?  core_alu_io_in1 :{ core_alu_io_in1 [0], core_alu_io_in1 [1], core_alu_io_in1 [2], core_alu_io_in1 [3], core_alu_io_in1 [4], core_alu__GEN_0 [18:15]|{ core_alu_io_in1 [7:6], core_alu_io_in1 [9:8]}&4'h5, core_alu__GEN_0 [14:7]| core_alu__GEN &8'h55, core_alu__GEN [1], core_alu__GEN_0 [5]| core_alu_io_in1 [18], core_alu_io_in1 [19], core_alu_io_in1 [20],{ core_alu__GEN_0 [2:0],1'h0}|{ core_alu_io_in1 [23:22], core_alu_io_in1 [25:24]}&4'h5, core_alu_io_in1 [25], core_alu_io_in1 [26], core_alu_io_in1 [27], core_alu_io_in1 [28], core_alu_io_in1 [29], core_alu_io_in1 [30], core_alu_io_in1 [31]}; 
    wire[32:0] core_alu__shout_r_T_5 =$signed($signed({ core_alu_io_fn [3]& core_alu_shin [31], core_alu_shin })>>> core_alu_shamt ); 
    wire[31:0] core_alu_shout_r = core_alu__shout_r_T_5 [31:0]; 
    wire[7:0] core_alu__GEN_1 ={{ core_alu_shout_r [11:8], core_alu_shout_r [15:14]}&6'h33,2'h0}|{ core_alu_shout_r [15:12], core_alu_shout_r [19:16]}&8'h33; 
    wire[18:0] core_alu__GEN_2 ={ core_alu_shout_r [5:4], core_alu_shout_r [7:6], core_alu_shout_r [9:8], core_alu__GEN_1 , core_alu_shout_r [19:18], core_alu_shout_r [21:20], core_alu_shout_r [23]}&19'h55555; 
    wire[31:0] core_alu_shout_l ={ core_alu_shout_r [0], core_alu_shout_r [1], core_alu_shout_r [2], core_alu_shout_r [3], core_alu_shout_r [4], core_alu__GEN_2 [18:15]|{ core_alu_shout_r [7:6], core_alu_shout_r [9:8]}&4'h5, core_alu__GEN_2 [14:7]| core_alu__GEN_1 &8'h55, core_alu__GEN_1 [1], core_alu__GEN_2 [5]| core_alu_shout_r [18], core_alu_shout_r [19], core_alu_shout_r [20],{ core_alu__GEN_2 [2:0],1'h0}|{ core_alu_shout_r [23:22], core_alu_shout_r [25:24]}&4'h5, core_alu_shout_r [25], core_alu_shout_r [26], core_alu_shout_r [27], core_alu_shout_r [28], core_alu_shout_r [29], core_alu_shout_r [30], core_alu_shout_r [31]}; 
    wire[31:0] core_alu_shout =( core_alu__shout_T | core_alu__shout_T_1  ?  core_alu_shout_r :32'h0)|( core_alu_io_fn ==4'h1 ?  core_alu_shout_l :32'h0); 
    wire core_alu_in2_not_zero =| core_alu_io_in2 ; 
    wire core_alu__logic_T_4 = core_alu_io_fn ==4'h6; 
    wire[31:0] core_alu_logic_0 =( core_alu_io_fn ==4'h4| core_alu__logic_T_4  ?  core_alu_in1_xor_in2 :32'h0)|( core_alu__logic_T_4 | core_alu_io_fn ==4'h7 ?  core_alu_io_in1 & core_alu_io_in2 :32'h0); 
    wire[31:0] core_alu_shift_logic ={31'h0, core_alu_io_fn >4'hB& core_alu_slt }| core_alu_logic_0 | core_alu_shout ; 
    wire[31:0] core_alu_out = core_alu_io_fn ==4'h0| core_alu_io_fn ==4'hA ?  core_alu__io_adder_out_T_3 : core_alu_shift_logic ; 
  assign  core_alu_io_out = core_alu_out ; 
  assign  core_alu_io_adder_out = core_alu__io_adder_out_T_3 ; 
  assign  core_alu_io_cmp_out = core_alu_io_fn [0]^( core_alu_io_fn [3] ?  core_alu_slt : core_alu_in1_xor_in2 ==32'h0);
    assign core_alu_io_fn = core_ex_ctrl_alu_fn;
    assign core_alu_io_in2 = core_ex_op2;
    assign core_alu_io_in1 = core_ex_op1;
    assign core__alu_io_out = core_alu_io_out;
    assign core_io_dmem_req_bits_addr = core_alu_io_adder_out;
    assign core__alu_io_cmp_out = core_alu_io_cmp_out;
      
    wire core_div_clock;
    wire core_div_reset;
    wire core_div_io_req_ready;
    wire core_div_io_req_valid;
    wire[3:0] core_div_io_req_bits_fn;
    wire core_div_io_req_bits_dw;
    wire[31:0] core_div_io_req_bits_in1;
    wire[31:0] core_div_io_req_bits_in2;
    wire[4:0] core_div_io_req_bits_tag;
    wire core_div_io_kill;
    wire core_div_io_resp_ready;
    wire core_div_io_resp_valid;
    wire[31:0] core_div_io_resp_bits_data;
    wire[4:0] core_div_io_resp_bits_tag;

    wire core_div_eOut =1'h0; reg[2:0] core_div_state ; reg[3:0] core_div_req_fn ; 
    reg core_div_req_dw ; reg[31:0] core_div_req_in1 ; reg[31:0] core_div_req_in2 ; reg[4:0] core_div_req_tag ; reg[5:0] core_div_count ; 
    reg core_div_neg_out ; 
    reg core_div_isHi ; 
    reg core_div_resHi ; reg[32:0] core_div_divisor ; 
    wire[32:0] core_div_mpcand = core_div_divisor ; reg[65:0] core_div_remainder ; 
    wire[2:0] core_div_decoded_plaInput ; 
    wire[2:0] core_div_decoded_invInputs =~ core_div_decoded_plaInput ; 
    wire[3:0] core_div_decoded_invMatrixOutputs ; 
    wire core_div_decoded_andMatrixInput_0 = core_div_decoded_invInputs [0]; 
    wire core_div_decoded_andMatrixInput_0_5 = core_div_decoded_invInputs [0]; 
    wire core_div_decoded_andMatrixInput_0_1 = core_div_decoded_invInputs [2]; 
    wire core_div_decoded_andMatrixInput_1 = core_div_decoded_invInputs [2]; 
    wire core_div_decoded_andMatrixInput_1_1 = core_div_decoded_invInputs [2]; 
    wire core_div_decoded_andMatrixInput_0_2 = core_div_decoded_invInputs [1]; 
    wire[1:0] core_div__decoded_T_2 ={ core_div_decoded_andMatrixInput_0_2 , core_div_decoded_andMatrixInput_1 }; 
    wire core_div_decoded_andMatrixInput_0_3 = core_div_decoded_plaInput [0]; 
    wire core_div_decoded_andMatrixInput_0_4 = core_div_decoded_plaInput [1]; 
    wire core_div_decoded_andMatrixInput_1_2 = core_div_decoded_plaInput [2]; 
    wire[1:0] core_div_decoded_orMatrixOutputs_lo ={|{ core_div_decoded_andMatrixInput_0 ,& core_div__decoded_T_2 },|{& core_div__decoded_T_2 ,&{ core_div_decoded_andMatrixInput_0_5 , core_div_decoded_andMatrixInput_1_2 }}}; 
    wire[1:0] core_div_decoded_orMatrixOutputs_hi ={ core_div_decoded_andMatrixInput_0_1 ,|{&{ core_div_decoded_andMatrixInput_0_3 , core_div_decoded_andMatrixInput_1_1 }, core_div_decoded_andMatrixInput_0_4 }}; 
    wire[3:0] core_div_decoded_orMatrixOutputs ={ core_div_decoded_orMatrixOutputs_hi , core_div_decoded_orMatrixOutputs_lo }; 
    wire[1:0] core_div_decoded_invMatrixOutputs_lo = core_div_decoded_orMatrixOutputs [1:0]; 
    wire[1:0] core_div_decoded_invMatrixOutputs_hi = core_div_decoded_orMatrixOutputs [3:2]; 
  assign  core_div_decoded_invMatrixOutputs ={ core_div_decoded_invMatrixOutputs_hi , core_div_decoded_invMatrixOutputs_lo }; 
    wire[3:0] core_div_decoded = core_div_decoded_invMatrixOutputs ; 
  assign  core_div_decoded_plaInput = core_div_io_req_bits_fn [2:0]; 
    wire core_div_cmdMul = core_div_decoded [3]; 
    wire core_div_cmdHi = core_div_decoded [2]; 
    wire core_div_lhsSigned = core_div_decoded [1]; 
    wire core_div_rhsSigned = core_div_decoded [0]; 
    wire core_div_lhs_sign = core_div_lhsSigned & core_div_io_req_bits_in1 [31]; 
    wire[15:0] core_div_hi = core_div_io_req_bits_in1 [31:16]; 
    wire[31:0] core_div_lhs_in ={ core_div_hi , core_div_io_req_bits_in1 [15:0]}; 
    wire core_div_rhs_sign = core_div_rhsSigned & core_div_io_req_bits_in2 [31]; 
    wire[15:0] core_div_hi_1 = core_div_io_req_bits_in2 [31:16]; 
    wire[31:0] core_div_rhs_in ={ core_div_hi_1 , core_div_io_req_bits_in2 [15:0]}; 
    wire[32:0] core_div_subtractor = core_div_remainder [64:32]- core_div_divisor ; 
    wire[31:0] core_div_result = core_div_resHi  ?  core_div_remainder [64:33]: core_div_remainder [31:0]; 
    wire[31:0] core_div_negated_remainder =32'h0- core_div_result ; 
    wire[64:0] core_div_mulReg ={ core_div_remainder [65:33], core_div_remainder [31:0]}; 
    wire core_div_mplierSign = core_div_remainder [32]; 
    wire[31:0] core_div_mplier = core_div_mulReg [31:0]; 
    wire[32:0] core_div_accum = core_div_mulReg [64:32]; 
    wire[41:0] core_div_prod ={{34{ core_div_mplierSign }}, core_div_mplier [7:0]}*{{9{ core_div_mpcand [32]}}, core_div_mpcand }+{{9{ core_div_accum [32]}}, core_div_accum }; 
    wire[41:0] core_div_nextMulReg_hi = core_div_prod ; 
    wire[65:0] core_div_nextMulReg ={ core_div_nextMulReg_hi , core_div_mplier [31:8]}; 
    wire core_div_nextMplierSign = core_div_count ==6'h2& core_div_neg_out ; 
    wire[32:0] core_div__eOutMask_T_2 =$signed(33'sh100000000>>>{28'h0, core_div_count [1:0],3'h0}); 
    wire[31:0] core_div_eOutMask = core_div__eOutMask_T_2 [31:0]; 
    wire[64:0] core_div_eOutRes = core_div_mulReg >>5'h0-{ core_div_count [1:0],3'h0}; 
    wire[64:0] core_div_nextMulReg1 = core_div_nextMulReg [64:0]; 
    wire[33:0] core_div_remainder_hi ={ core_div_nextMulReg1 [64:32], core_div_nextMplierSign }; 
    wire core_div_unrolls_less = core_div_subtractor [32]; 
    wire[63:0] core_div_unrolls_hi ={ core_div_unrolls_less  ?  core_div_remainder [63:32]: core_div_subtractor [31:0], core_div_remainder [31:0]}; 
    wire[64:0] core_div_unrolls_0 ={ core_div_unrolls_hi ,~ core_div_unrolls_less }; 
    wire core_div_divby0 = core_div_count ==6'h0&~ core_div_unrolls_less ; 
    wire core_div_outMul =~( core_div_state [0]); 
    wire[15:0] core_div_hiOut = core_div_result [31:16]; 
    wire[15:0] core_div_loOut = core_div_result [15:0]; 
    wire core_div__io_resp_valid_output = core_div_state ==3'h6|(& core_div_state ); 
    wire core_div__io_req_ready_output = core_div_state ==3'h0; 
    wire core_div__GEN = core_div_state ==3'h1; 
    wire core_div__GEN_0 = core_div_state ==3'h5; 
    wire core_div__GEN_1 = core_div_state ==3'h2; 
    wire core_div__GEN_2 = core_div__GEN_1 & core_div_count ==6'h3; 
    wire core_div__GEN_3 = core_div_state ==3'h3; 
    wire core_div__GEN_4 = core_div_count ==6'h20; 
    wire core_div__GEN_5 = core_div__io_req_ready_output & core_div_io_req_valid ; 
  always @( posedge  core_div_clock )
         begin 
             if ( core_div_reset ) 
                 core_div_state  <=3'h0;
              else 
                 if ( core_div__GEN_5 ) 
                     core_div_state  <= core_div_cmdMul  ? 3'h2:{1'h0,~( core_div_lhs_sign | core_div_rhs_sign ),1'h1};
                  else 
                     if ( core_div_io_resp_ready & core_div__io_resp_valid_output | core_div_io_kill ) 
                         core_div_state  <=3'h0;
                      else 
                         if ( core_div__GEN_3 & core_div__GEN_4 ) 
                             core_div_state  <={1'h1,~ core_div_neg_out ,1'h1};
                          else 
                             if ( core_div__GEN_2 ) 
                                 core_div_state  <=3'h6;
                              else 
                                 if ( core_div__GEN_0 ) 
                                     core_div_state  <=3'h7;
                                  else 
                                     if ( core_div__GEN ) 
                                         core_div_state  <=3'h3;
             if ( core_div__GEN_5 )
                 begin  
                     core_div_req_fn  <= core_div_io_req_bits_fn ; 
                     core_div_req_dw  <= core_div_io_req_bits_dw ; 
                     core_div_req_in1  <= core_div_io_req_bits_in1 ; 
                     core_div_req_in2  <= core_div_io_req_bits_in2 ; 
                     core_div_req_tag  <= core_div_io_req_bits_tag ; 
                     core_div_count  <=6'h0; 
                     core_div_neg_out  <= core_div_cmdHi  ?  core_div_lhs_sign : core_div_lhs_sign != core_div_rhs_sign ; 
                     core_div_isHi  <= core_div_cmdHi ; 
                     core_div_divisor  <={ core_div_rhs_sign , core_div_rhs_in }; 
                     core_div_remainder  <={34'h0, core_div_lhs_in };
                 end 
              else 
                 begin 
                     if ( core_div__GEN_3 )
                         begin  
                             core_div_count  <= core_div_count +6'h1; 
                             core_div_remainder  <={1'h0, core_div_unrolls_0 };
                         end 
                      else 
                         if ( core_div__GEN_1 )
                             begin  
                                 core_div_count  <= core_div_count +6'h1; 
                                 core_div_remainder  <={ core_div_remainder_hi , core_div_nextMulReg1 [31:0]};
                             end 
                          else 
                             if ( core_div__GEN_0 | core_div__GEN & core_div_remainder [31]) 
                                 core_div_remainder  <={34'h0, core_div_negated_remainder }; 
                     core_div_neg_out  <=~( core_div__GEN_3 & core_div_divby0 &~ core_div_isHi )& core_div_neg_out ;
                     if ( core_div__GEN & core_div_divisor [31]) 
                         core_div_divisor  <= core_div_subtractor ;
                 end  
             core_div_resHi  <=~ core_div__GEN_5 &( core_div__GEN_3 & core_div__GEN_4 | core_div__GEN_2  ?  core_div_isHi :~ core_div__GEN_0 & core_div_resHi );
         end
  assign  core_div_io_req_ready = core_div__io_req_ready_output ; 
  assign  core_div_io_resp_valid = core_div__io_resp_valid_output ; 
  assign  core_div_io_resp_bits_data ={ core_div_hiOut , core_div_loOut }; 
  assign  core_div_io_resp_bits_tag = core_div_req_tag ;
    assign core_div_clock = core_clock;
    assign core_div_reset = core_reset;
    assign core__div_io_req_ready = core_div_io_req_ready;
    assign core_div_io_req_valid = core__div_io_req_valid_T;
    assign core_div_io_req_bits_fn = core_ex_ctrl_alu_fn;
    assign core_div_io_req_bits_dw = core_ex_ctrl_alu_dw;
    assign core_div_io_req_bits_in1 = core_ex_rs_0;
    assign core_div_io_req_bits_in2 = core_ex_rs_1;
    assign core_div_io_req_bits_tag = core_ex_waddr;
    assign core_div_io_kill = core_killm_common&core_div_io_kill_REG;
    assign core_div_io_resp_ready = core__GEN;
    assign core__div_io_resp_valid = core_div_io_resp_valid;
    assign core_ll_wdata = core_div_io_resp_bits_data;
    assign core__div_io_resp_bits_tag = core_div_io_resp_bits_tag;
      
    wire core_PlusArgTimeout_clock;
    wire core_PlusArgTimeout_reset;
    wire[31:0] core_PlusArgTimeout_io_count;

    wire[31:0] core_PlusArgTimeout__plusarg_reader_out ; 
  always @( posedge  core_PlusArgTimeout_clock )
         begin 
             if ((| core_PlusArgTimeout__plusarg_reader_out )&~ core_PlusArgTimeout_reset & core_PlusArgTimeout_io_count >= core_PlusArgTimeout__plusarg_reader_out )
                 begin 
                     if (1)$error("Assertion failed: Timeout exceeded: Kill the emulation after INT rdtime cycles. Off if 0.\n    at PlusArg.scala:64 assert (io.count < max, s\"Timeout exceeded: $docstring\")\n");
                     if (1)$fatal;
                 end 
         end
    plusarg_reader  #(. core_PlusArgTimeout_DEFAULT (0),. core_PlusArgTimeout_FORMAT ("max_core_cycles=%d"),. core_PlusArgTimeout_WIDTH (32)) core_PlusArgTimeout_plusarg_reader (. out ( core_PlusArgTimeout__plusarg_reader_out ));
    assign core_PlusArgTimeout_clock = core_clock;
    assign core_PlusArgTimeout_reset = core_reset;
    assign core_PlusArgTimeout_io_count = core__csr_io_time;
     
  assign  core_io_imem_might_request = core_imem_might_request_reg ; 
  assign  core_io_imem_req_valid = core_take_pc_mem_wb ; 
  assign  core_io_imem_req_bits_pc = core_wb_xcpt | core__csr_io_eret  ?  core__csr_io_evec : core_replay_wb  ?  core_wb_reg_pc : core_mem_npc ; 
  assign  core_io_imem_req_bits_speculative =~ core_take_pc_wb ; 
  assign  core_io_imem_sfence_valid = core__io_imem_sfence_valid_output ; 
  assign  core_io_imem_btb_update_valid = core_mem_reg_valid &~ core_take_pc_wb & core_mem_wrong_npc &(~ core_mem_cfi | core_mem_cfi_taken ); 
  assign  core_io_imem_bht_update_valid = core_mem_reg_valid &~ core_take_pc_wb ; 
  assign  core_io_imem_flush_icache = core_wb_reg_valid & core_wb_ctrl_fence_i &~ core_io_dmem_s2_nack ; 
  assign  core_io_imem_progress = core_io_imem_progress_REG ; 
  assign  core_io_dmem_req_valid = core__io_dmem_req_valid_output ; 
  assign  core_io_dmem_req_bits_tag ={1'h0, core_ex_dcache_tag }; 
  assign  core_io_dmem_req_bits_cmd = core_ex_ctrl_mem_cmd ; 
  assign  core_io_dmem_req_bits_size = core_ex_reg_mem_size ; 
  assign  core_io_dmem_req_bits_signed =~( core_ex_reg_inst [14]); 
  assign  core_io_dmem_req_bits_dv = core__csr_io_status_dv ; 
  assign  core_io_dmem_s1_kill = core_killm_common | core_mem_ldst_xcpt ; 
  assign  core_io_dmem_s1_data_data = core_mem_reg_rs2 ; 
  assign  core_io_ptw_sfence_valid = core__io_imem_sfence_valid_output ; 
  assign  core_io_ptw_sfence_bits_rs1 = core_wb_reg_mem_size [0]; 
  assign  core_io_ptw_status_debug = core__csr_io_status_debug ; 
  assign  core_io_ptw_customCSRs_csrs_0_value = core__csr_io_customCSRs_0_value ; 
  assign  core_io_trace_insns_0_valid = core__csr_io_trace_0_valid ; 
  assign  core_io_trace_insns_0_iaddr = core__csr_io_trace_0_iaddr ; 
  assign  core_io_trace_insns_0_insn = core__csr_io_trace_0_insn ; 
  assign  core_io_trace_insns_0_priv = core__csr_io_trace_0_priv ; 
  assign  core_io_trace_insns_0_exception = core__csr_io_trace_0_exception ; 
  assign  core_io_trace_time ={32'h0, core__csr_io_time }; 
  assign  core_io_bpwatch_0_valid_0 = core_wb_reg_wphit_0 ; 
  assign  core_io_bpwatch_0_action ={2'h0, core__csr_io_bp_0_control_action };
    assign core_clock = clock;
    assign core_reset = reset;
    assign core_io_hartid = hartIdSinkNodeIn;
    assign core_io_interrupts_debug = intSinkNodeIn_0;
    assign core_io_interrupts_mtip = intSinkNodeIn_2;
    assign core_io_interrupts_msip = intSinkNodeIn_1;
    assign core_io_interrupts_meip = intSinkNodeIn_3;
    assign _core_io_imem_might_request = core_io_imem_might_request;
    assign _core_io_imem_req_valid = core_io_imem_req_valid;
    assign _core_io_imem_req_bits_pc = core_io_imem_req_bits_pc;
    assign _core_io_imem_req_bits_speculative = core_io_imem_req_bits_speculative;
    assign _core_io_imem_sfence_valid = core_io_imem_sfence_valid;
    assign _core_io_imem_resp_ready = core_io_imem_resp_ready;
    assign core_io_imem_resp_valid = _frontend_io_cpu_resp_valid;
    assign core_io_imem_resp_bits_btb_cfiType = _frontend_io_cpu_resp_bits_btb_cfiType;
    assign core_io_imem_resp_bits_btb_taken = _frontend_io_cpu_resp_bits_btb_taken;
    assign core_io_imem_resp_bits_btb_mask = _frontend_io_cpu_resp_bits_btb_mask;
    assign core_io_imem_resp_bits_btb_bridx = _frontend_io_cpu_resp_bits_btb_bridx;
    assign core_io_imem_resp_bits_btb_target = _frontend_io_cpu_resp_bits_btb_target;
    assign core_io_imem_resp_bits_btb_entry = _frontend_io_cpu_resp_bits_btb_entry;
    assign core_io_imem_resp_bits_btb_bht_history = _frontend_io_cpu_resp_bits_btb_bht_history;
    assign core_io_imem_resp_bits_btb_bht_value = _frontend_io_cpu_resp_bits_btb_bht_value;
    assign core_io_imem_resp_bits_pc = _frontend_io_cpu_resp_bits_pc;
    assign core_io_imem_resp_bits_data = _frontend_io_cpu_resp_bits_data;
    assign core_io_imem_resp_bits_mask = _frontend_io_cpu_resp_bits_mask;
    assign core_io_imem_resp_bits_xcpt_pf_inst = _frontend_io_cpu_resp_bits_xcpt_pf_inst;
    assign core_io_imem_resp_bits_xcpt_gf_inst = _frontend_io_cpu_resp_bits_xcpt_gf_inst;
    assign core_io_imem_resp_bits_xcpt_ae_inst = _frontend_io_cpu_resp_bits_xcpt_ae_inst;
    assign core_io_imem_resp_bits_replay = _frontend_io_cpu_resp_bits_replay;
    assign core_io_imem_gpa_valid = _frontend_io_cpu_gpa_valid;
    assign core_io_imem_gpa_bits = _frontend_io_cpu_gpa_bits;
    assign _core_io_imem_btb_update_valid = core_io_imem_btb_update_valid;
    assign _core_io_imem_bht_update_valid = core_io_imem_bht_update_valid;
    assign _core_io_imem_flush_icache = core_io_imem_flush_icache;
    assign _core_io_imem_progress = core_io_imem_progress;
    assign core_io_dmem_req_ready = _dcacheArb_io_requestor_0_req_ready;
    assign _core_io_dmem_req_valid = core_io_dmem_req_valid;
    assign _core_io_dmem_req_bits_addr = core_io_dmem_req_bits_addr;
    assign _core_io_dmem_req_bits_tag = core_io_dmem_req_bits_tag;
    assign _core_io_dmem_req_bits_cmd = core_io_dmem_req_bits_cmd;
    assign _core_io_dmem_req_bits_size = core_io_dmem_req_bits_size;
    assign _core_io_dmem_req_bits_signed = core_io_dmem_req_bits_signed;
    assign _core_io_dmem_req_bits_dv = core_io_dmem_req_bits_dv;
    assign _core_io_dmem_s1_kill = core_io_dmem_s1_kill;
    assign _core_io_dmem_s1_data_data = core_io_dmem_s1_data_data;
    assign core_io_dmem_s2_nack = _dcacheArb_io_requestor_0_s2_nack;
    assign core_io_dmem_resp_valid = _dcacheArb_io_requestor_0_resp_valid;
    assign core_io_dmem_resp_bits_tag = _dcacheArb_io_requestor_0_resp_bits_tag;
    assign core_io_dmem_resp_bits_data = _dcacheArb_io_requestor_0_resp_bits_data;
    assign core_io_dmem_resp_bits_replay = _dcacheArb_io_requestor_0_resp_bits_replay;
    assign core_io_dmem_resp_bits_has_data = _dcacheArb_io_requestor_0_resp_bits_has_data;
    assign core_io_dmem_resp_bits_data_word_bypass = _dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
    assign core_io_dmem_replay_next = _dcacheArb_io_requestor_0_replay_next;
    assign core_io_dmem_s2_xcpt_ma_ld = _dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
    assign core_io_dmem_s2_xcpt_ma_st = _dcacheArb_io_requestor_0_s2_xcpt_ma_st;
    assign core_io_dmem_s2_xcpt_pf_ld = _dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
    assign core_io_dmem_s2_xcpt_pf_st = _dcacheArb_io_requestor_0_s2_xcpt_pf_st;
    assign core_io_dmem_s2_xcpt_ae_ld = _dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
    assign core_io_dmem_s2_xcpt_ae_st = _dcacheArb_io_requestor_0_s2_xcpt_ae_st;
    assign core_io_dmem_ordered = _dcacheArb_io_requestor_0_ordered;
    assign core_io_dmem_perf_grant = _dcacheArb_io_requestor_0_perf_grant;
    assign _core_io_ptw_sfence_valid = core_io_ptw_sfence_valid;
    assign _core_io_ptw_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1;
    assign _core_io_ptw_status_debug = core_io_ptw_status_debug;
    assign _core_io_ptw_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l;
    assign _core_io_ptw_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a;
    assign _core_io_ptw_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x;
    assign _core_io_ptw_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w;
    assign _core_io_ptw_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r;
    assign _core_io_ptw_pmp_0_addr = core_io_ptw_pmp_0_addr;
    assign _core_io_ptw_pmp_0_mask = core_io_ptw_pmp_0_mask;
    assign _core_io_ptw_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l;
    assign _core_io_ptw_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a;
    assign _core_io_ptw_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x;
    assign _core_io_ptw_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w;
    assign _core_io_ptw_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r;
    assign _core_io_ptw_pmp_1_addr = core_io_ptw_pmp_1_addr;
    assign _core_io_ptw_pmp_1_mask = core_io_ptw_pmp_1_mask;
    assign _core_io_ptw_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l;
    assign _core_io_ptw_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a;
    assign _core_io_ptw_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x;
    assign _core_io_ptw_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w;
    assign _core_io_ptw_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r;
    assign _core_io_ptw_pmp_2_addr = core_io_ptw_pmp_2_addr;
    assign _core_io_ptw_pmp_2_mask = core_io_ptw_pmp_2_mask;
    assign _core_io_ptw_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l;
    assign _core_io_ptw_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a;
    assign _core_io_ptw_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x;
    assign _core_io_ptw_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w;
    assign _core_io_ptw_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r;
    assign _core_io_ptw_pmp_3_addr = core_io_ptw_pmp_3_addr;
    assign _core_io_ptw_pmp_3_mask = core_io_ptw_pmp_3_mask;
    assign _core_io_ptw_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l;
    assign _core_io_ptw_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a;
    assign _core_io_ptw_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x;
    assign _core_io_ptw_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w;
    assign _core_io_ptw_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r;
    assign _core_io_ptw_pmp_4_addr = core_io_ptw_pmp_4_addr;
    assign _core_io_ptw_pmp_4_mask = core_io_ptw_pmp_4_mask;
    assign _core_io_ptw_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l;
    assign _core_io_ptw_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a;
    assign _core_io_ptw_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x;
    assign _core_io_ptw_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w;
    assign _core_io_ptw_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r;
    assign _core_io_ptw_pmp_5_addr = core_io_ptw_pmp_5_addr;
    assign _core_io_ptw_pmp_5_mask = core_io_ptw_pmp_5_mask;
    assign _core_io_ptw_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l;
    assign _core_io_ptw_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a;
    assign _core_io_ptw_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x;
    assign _core_io_ptw_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w;
    assign _core_io_ptw_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r;
    assign _core_io_ptw_pmp_6_addr = core_io_ptw_pmp_6_addr;
    assign _core_io_ptw_pmp_6_mask = core_io_ptw_pmp_6_mask;
    assign _core_io_ptw_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l;
    assign _core_io_ptw_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a;
    assign _core_io_ptw_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x;
    assign _core_io_ptw_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w;
    assign _core_io_ptw_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r;
    assign _core_io_ptw_pmp_7_addr = core_io_ptw_pmp_7_addr;
    assign _core_io_ptw_pmp_7_mask = core_io_ptw_pmp_7_mask;
    assign _core_io_ptw_customCSRs_csrs_0_value = core_io_ptw_customCSRs_csrs_0_value;
    assign traceSourceNodeOut_insns_0_valid = core_io_trace_insns_0_valid;
    assign traceSourceNodeOut_insns_0_iaddr = core_io_trace_insns_0_iaddr;
    assign traceSourceNodeOut_insns_0_insn = core_io_trace_insns_0_insn;
    assign traceSourceNodeOut_insns_0_priv = core_io_trace_insns_0_priv;
    assign traceSourceNodeOut_insns_0_exception = core_io_trace_insns_0_exception;
    assign traceSourceNodeOut_insns_0_interrupt = core_io_trace_insns_0_interrupt;
    assign traceSourceNodeOut_insns_0_cause = core_io_trace_insns_0_cause;
    assign traceSourceNodeOut_insns_0_tval = core_io_trace_insns_0_tval;
    assign traceSourceNodeOut_time = core_io_trace_time;
    assign bpwatchSourceNodeOut_0_valid_0 = core_io_bpwatch_0_valid_0;
    assign bpwatchSourceNodeOut_0_action = core_io_bpwatch_0_action;
    assign _core_io_wfi = core_io_wfi;
    
  assign auto_buffer_in_a_ready = buffer_1_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign auto_buffer_in_d_valid = buffer_1_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign auto_buffer_in_d_bits_opcode = buffer_1_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign auto_buffer_in_d_bits_size = buffer_1_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign auto_buffer_in_d_bits_source = buffer_1_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign auto_buffer_in_d_bits_data = buffer_1_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign auto_buffer_out_a_valid = buffer_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_opcode = buffer_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_param = buffer_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_size = buffer_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_source = buffer_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_address = buffer_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_mask = buffer_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_a_bits_data = buffer_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_buffer_out_d_ready = buffer_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_valid = broadcast_3_nodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_iaddr = broadcast_3_nodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_insn = broadcast_3_nodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_priv = broadcast_3_nodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_exception = broadcast_3_nodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_interrupt = broadcast_3_nodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_cause = broadcast_3_nodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_insns_0_tval = broadcast_3_nodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_broadcast_out_time = broadcast_3_nodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_wfi_out_0 = wfiNodeOut_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
endmodule